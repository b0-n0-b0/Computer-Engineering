library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity ddfs_lut_4096_6bit is
  port (
    address  : in  std_logic_vector(11 downto 0);
    ddfs_out : out std_logic_vector(5 downto 0)
  );
end entity;

architecture rtl of ddfs_lut_4096_6bit is

  type LUT_t is array (natural range 0 to 4095) of integer;
  constant LUT: LUT_t := (
    0 => 0,
    1 => 0,
    2 => 0,
    3 => 0,
    4 => 0,
    5 => 0,
    6 => 0,
    7 => 0,
    8 => 0,
    9 => 0,
    10 => 0,
    11 => 1,
    12 => 1,
    13 => 1,
    14 => 1,
    15 => 1,
    16 => 1,
    17 => 1,
    18 => 1,
    19 => 1,
    20 => 1,
    21 => 1,
    22 => 1,
    23 => 1,
    24 => 1,
    25 => 1,
    26 => 1,
    27 => 1,
    28 => 1,
    29 => 1,
    30 => 1,
    31 => 1,
    32 => 2,
    33 => 2,
    34 => 2,
    35 => 2,
    36 => 2,
    37 => 2,
    38 => 2,
    39 => 2,
    40 => 2,
    41 => 2,
    42 => 2,
    43 => 2,
    44 => 2,
    45 => 2,
    46 => 2,
    47 => 2,
    48 => 2,
    49 => 2,
    50 => 2,
    51 => 2,
    52 => 2,
    53 => 3,
    54 => 3,
    55 => 3,
    56 => 3,
    57 => 3,
    58 => 3,
    59 => 3,
    60 => 3,
    61 => 3,
    62 => 3,
    63 => 3,
    64 => 3,
    65 => 3,
    66 => 3,
    67 => 3,
    68 => 3,
    69 => 3,
    70 => 3,
    71 => 3,
    72 => 3,
    73 => 3,
    74 => 4,
    75 => 4,
    76 => 4,
    77 => 4,
    78 => 4,
    79 => 4,
    80 => 4,
    81 => 4,
    82 => 4,
    83 => 4,
    84 => 4,
    85 => 4,
    86 => 4,
    87 => 4,
    88 => 4,
    89 => 4,
    90 => 4,
    91 => 4,
    92 => 4,
    93 => 4,
    94 => 4,
    95 => 5,
    96 => 5,
    97 => 5,
    98 => 5,
    99 => 5,
    100 => 5,
    101 => 5,
    102 => 5,
    103 => 5,
    104 => 5,
    105 => 5,
    106 => 5,
    107 => 5,
    108 => 5,
    109 => 5,
    110 => 5,
    111 => 5,
    112 => 5,
    113 => 5,
    114 => 5,
    115 => 5,
    116 => 5,
    117 => 6,
    118 => 6,
    119 => 6,
    120 => 6,
    121 => 6,
    122 => 6,
    123 => 6,
    124 => 6,
    125 => 6,
    126 => 6,
    127 => 6,
    128 => 6,
    129 => 6,
    130 => 6,
    131 => 6,
    132 => 6,
    133 => 6,
    134 => 6,
    135 => 6,
    136 => 6,
    137 => 6,
    138 => 7,
    139 => 7,
    140 => 7,
    141 => 7,
    142 => 7,
    143 => 7,
    144 => 7,
    145 => 7,
    146 => 7,
    147 => 7,
    148 => 7,
    149 => 7,
    150 => 7,
    151 => 7,
    152 => 7,
    153 => 7,
    154 => 7,
    155 => 7,
    156 => 7,
    157 => 7,
    158 => 7,
    159 => 7,
    160 => 8,
    161 => 8,
    162 => 8,
    163 => 8,
    164 => 8,
    165 => 8,
    166 => 8,
    167 => 8,
    168 => 8,
    169 => 8,
    170 => 8,
    171 => 8,
    172 => 8,
    173 => 8,
    174 => 8,
    175 => 8,
    176 => 8,
    177 => 8,
    178 => 8,
    179 => 8,
    180 => 8,
    181 => 8,
    182 => 9,
    183 => 9,
    184 => 9,
    185 => 9,
    186 => 9,
    187 => 9,
    188 => 9,
    189 => 9,
    190 => 9,
    191 => 9,
    192 => 9,
    193 => 9,
    194 => 9,
    195 => 9,
    196 => 9,
    197 => 9,
    198 => 9,
    199 => 9,
    200 => 9,
    201 => 9,
    202 => 9,
    203 => 9,
    204 => 10,
    205 => 10,
    206 => 10,
    207 => 10,
    208 => 10,
    209 => 10,
    210 => 10,
    211 => 10,
    212 => 10,
    213 => 10,
    214 => 10,
    215 => 10,
    216 => 10,
    217 => 10,
    218 => 10,
    219 => 10,
    220 => 10,
    221 => 10,
    222 => 10,
    223 => 10,
    224 => 10,
    225 => 10,
    226 => 11,
    227 => 11,
    228 => 11,
    229 => 11,
    230 => 11,
    231 => 11,
    232 => 11,
    233 => 11,
    234 => 11,
    235 => 11,
    236 => 11,
    237 => 11,
    238 => 11,
    239 => 11,
    240 => 11,
    241 => 11,
    242 => 11,
    243 => 11,
    244 => 11,
    245 => 11,
    246 => 11,
    247 => 11,
    248 => 12,
    249 => 12,
    250 => 12,
    251 => 12,
    252 => 12,
    253 => 12,
    254 => 12,
    255 => 12,
    256 => 12,
    257 => 12,
    258 => 12,
    259 => 12,
    260 => 12,
    261 => 12,
    262 => 12,
    263 => 12,
    264 => 12,
    265 => 12,
    266 => 12,
    267 => 12,
    268 => 12,
    269 => 12,
    270 => 12,
    271 => 13,
    272 => 13,
    273 => 13,
    274 => 13,
    275 => 13,
    276 => 13,
    277 => 13,
    278 => 13,
    279 => 13,
    280 => 13,
    281 => 13,
    282 => 13,
    283 => 13,
    284 => 13,
    285 => 13,
    286 => 13,
    287 => 13,
    288 => 13,
    289 => 13,
    290 => 13,
    291 => 13,
    292 => 13,
    293 => 13,
    294 => 14,
    295 => 14,
    296 => 14,
    297 => 14,
    298 => 14,
    299 => 14,
    300 => 14,
    301 => 14,
    302 => 14,
    303 => 14,
    304 => 14,
    305 => 14,
    306 => 14,
    307 => 14,
    308 => 14,
    309 => 14,
    310 => 14,
    311 => 14,
    312 => 14,
    313 => 14,
    314 => 14,
    315 => 14,
    316 => 14,
    317 => 14,
    318 => 15,
    319 => 15,
    320 => 15,
    321 => 15,
    322 => 15,
    323 => 15,
    324 => 15,
    325 => 15,
    326 => 15,
    327 => 15,
    328 => 15,
    329 => 15,
    330 => 15,
    331 => 15,
    332 => 15,
    333 => 15,
    334 => 15,
    335 => 15,
    336 => 15,
    337 => 15,
    338 => 15,
    339 => 15,
    340 => 15,
    341 => 15,
    342 => 16,
    343 => 16,
    344 => 16,
    345 => 16,
    346 => 16,
    347 => 16,
    348 => 16,
    349 => 16,
    350 => 16,
    351 => 16,
    352 => 16,
    353 => 16,
    354 => 16,
    355 => 16,
    356 => 16,
    357 => 16,
    358 => 16,
    359 => 16,
    360 => 16,
    361 => 16,
    362 => 16,
    363 => 16,
    364 => 16,
    365 => 16,
    366 => 17,
    367 => 17,
    368 => 17,
    369 => 17,
    370 => 17,
    371 => 17,
    372 => 17,
    373 => 17,
    374 => 17,
    375 => 17,
    376 => 17,
    377 => 17,
    378 => 17,
    379 => 17,
    380 => 17,
    381 => 17,
    382 => 17,
    383 => 17,
    384 => 17,
    385 => 17,
    386 => 17,
    387 => 17,
    388 => 17,
    389 => 17,
    390 => 17,
    391 => 17,
    392 => 18,
    393 => 18,
    394 => 18,
    395 => 18,
    396 => 18,
    397 => 18,
    398 => 18,
    399 => 18,
    400 => 18,
    401 => 18,
    402 => 18,
    403 => 18,
    404 => 18,
    405 => 18,
    406 => 18,
    407 => 18,
    408 => 18,
    409 => 18,
    410 => 18,
    411 => 18,
    412 => 18,
    413 => 18,
    414 => 18,
    415 => 18,
    416 => 18,
    417 => 19,
    418 => 19,
    419 => 19,
    420 => 19,
    421 => 19,
    422 => 19,
    423 => 19,
    424 => 19,
    425 => 19,
    426 => 19,
    427 => 19,
    428 => 19,
    429 => 19,
    430 => 19,
    431 => 19,
    432 => 19,
    433 => 19,
    434 => 19,
    435 => 19,
    436 => 19,
    437 => 19,
    438 => 19,
    439 => 19,
    440 => 19,
    441 => 19,
    442 => 19,
    443 => 19,
    444 => 20,
    445 => 20,
    446 => 20,
    447 => 20,
    448 => 20,
    449 => 20,
    450 => 20,
    451 => 20,
    452 => 20,
    453 => 20,
    454 => 20,
    455 => 20,
    456 => 20,
    457 => 20,
    458 => 20,
    459 => 20,
    460 => 20,
    461 => 20,
    462 => 20,
    463 => 20,
    464 => 20,
    465 => 20,
    466 => 20,
    467 => 20,
    468 => 20,
    469 => 20,
    470 => 20,
    471 => 20,
    472 => 21,
    473 => 21,
    474 => 21,
    475 => 21,
    476 => 21,
    477 => 21,
    478 => 21,
    479 => 21,
    480 => 21,
    481 => 21,
    482 => 21,
    483 => 21,
    484 => 21,
    485 => 21,
    486 => 21,
    487 => 21,
    488 => 21,
    489 => 21,
    490 => 21,
    491 => 21,
    492 => 21,
    493 => 21,
    494 => 21,
    495 => 21,
    496 => 21,
    497 => 21,
    498 => 21,
    499 => 21,
    500 => 22,
    501 => 22,
    502 => 22,
    503 => 22,
    504 => 22,
    505 => 22,
    506 => 22,
    507 => 22,
    508 => 22,
    509 => 22,
    510 => 22,
    511 => 22,
    512 => 22,
    513 => 22,
    514 => 22,
    515 => 22,
    516 => 22,
    517 => 22,
    518 => 22,
    519 => 22,
    520 => 22,
    521 => 22,
    522 => 22,
    523 => 22,
    524 => 22,
    525 => 22,
    526 => 22,
    527 => 22,
    528 => 22,
    529 => 22,
    530 => 23,
    531 => 23,
    532 => 23,
    533 => 23,
    534 => 23,
    535 => 23,
    536 => 23,
    537 => 23,
    538 => 23,
    539 => 23,
    540 => 23,
    541 => 23,
    542 => 23,
    543 => 23,
    544 => 23,
    545 => 23,
    546 => 23,
    547 => 23,
    548 => 23,
    549 => 23,
    550 => 23,
    551 => 23,
    552 => 23,
    553 => 23,
    554 => 23,
    555 => 23,
    556 => 23,
    557 => 23,
    558 => 23,
    559 => 23,
    560 => 23,
    561 => 24,
    562 => 24,
    563 => 24,
    564 => 24,
    565 => 24,
    566 => 24,
    567 => 24,
    568 => 24,
    569 => 24,
    570 => 24,
    571 => 24,
    572 => 24,
    573 => 24,
    574 => 24,
    575 => 24,
    576 => 24,
    577 => 24,
    578 => 24,
    579 => 24,
    580 => 24,
    581 => 24,
    582 => 24,
    583 => 24,
    584 => 24,
    585 => 24,
    586 => 24,
    587 => 24,
    588 => 24,
    589 => 24,
    590 => 24,
    591 => 24,
    592 => 24,
    593 => 24,
    594 => 24,
    595 => 25,
    596 => 25,
    597 => 25,
    598 => 25,
    599 => 25,
    600 => 25,
    601 => 25,
    602 => 25,
    603 => 25,
    604 => 25,
    605 => 25,
    606 => 25,
    607 => 25,
    608 => 25,
    609 => 25,
    610 => 25,
    611 => 25,
    612 => 25,
    613 => 25,
    614 => 25,
    615 => 25,
    616 => 25,
    617 => 25,
    618 => 25,
    619 => 25,
    620 => 25,
    621 => 25,
    622 => 25,
    623 => 25,
    624 => 25,
    625 => 25,
    626 => 25,
    627 => 25,
    628 => 25,
    629 => 25,
    630 => 26,
    631 => 26,
    632 => 26,
    633 => 26,
    634 => 26,
    635 => 26,
    636 => 26,
    637 => 26,
    638 => 26,
    639 => 26,
    640 => 26,
    641 => 26,
    642 => 26,
    643 => 26,
    644 => 26,
    645 => 26,
    646 => 26,
    647 => 26,
    648 => 26,
    649 => 26,
    650 => 26,
    651 => 26,
    652 => 26,
    653 => 26,
    654 => 26,
    655 => 26,
    656 => 26,
    657 => 26,
    658 => 26,
    659 => 26,
    660 => 26,
    661 => 26,
    662 => 26,
    663 => 26,
    664 => 26,
    665 => 26,
    666 => 26,
    667 => 26,
    668 => 26,
    669 => 27,
    670 => 27,
    671 => 27,
    672 => 27,
    673 => 27,
    674 => 27,
    675 => 27,
    676 => 27,
    677 => 27,
    678 => 27,
    679 => 27,
    680 => 27,
    681 => 27,
    682 => 27,
    683 => 27,
    684 => 27,
    685 => 27,
    686 => 27,
    687 => 27,
    688 => 27,
    689 => 27,
    690 => 27,
    691 => 27,
    692 => 27,
    693 => 27,
    694 => 27,
    695 => 27,
    696 => 27,
    697 => 27,
    698 => 27,
    699 => 27,
    700 => 27,
    701 => 27,
    702 => 27,
    703 => 27,
    704 => 27,
    705 => 27,
    706 => 27,
    707 => 27,
    708 => 27,
    709 => 27,
    710 => 27,
    711 => 27,
    712 => 28,
    713 => 28,
    714 => 28,
    715 => 28,
    716 => 28,
    717 => 28,
    718 => 28,
    719 => 28,
    720 => 28,
    721 => 28,
    722 => 28,
    723 => 28,
    724 => 28,
    725 => 28,
    726 => 28,
    727 => 28,
    728 => 28,
    729 => 28,
    730 => 28,
    731 => 28,
    732 => 28,
    733 => 28,
    734 => 28,
    735 => 28,
    736 => 28,
    737 => 28,
    738 => 28,
    739 => 28,
    740 => 28,
    741 => 28,
    742 => 28,
    743 => 28,
    744 => 28,
    745 => 28,
    746 => 28,
    747 => 28,
    748 => 28,
    749 => 28,
    750 => 28,
    751 => 28,
    752 => 28,
    753 => 28,
    754 => 28,
    755 => 28,
    756 => 28,
    757 => 28,
    758 => 28,
    759 => 28,
    760 => 28,
    761 => 29,
    762 => 29,
    763 => 29,
    764 => 29,
    765 => 29,
    766 => 29,
    767 => 29,
    768 => 29,
    769 => 29,
    770 => 29,
    771 => 29,
    772 => 29,
    773 => 29,
    774 => 29,
    775 => 29,
    776 => 29,
    777 => 29,
    778 => 29,
    779 => 29,
    780 => 29,
    781 => 29,
    782 => 29,
    783 => 29,
    784 => 29,
    785 => 29,
    786 => 29,
    787 => 29,
    788 => 29,
    789 => 29,
    790 => 29,
    791 => 29,
    792 => 29,
    793 => 29,
    794 => 29,
    795 => 29,
    796 => 29,
    797 => 29,
    798 => 29,
    799 => 29,
    800 => 29,
    801 => 29,
    802 => 29,
    803 => 29,
    804 => 29,
    805 => 29,
    806 => 29,
    807 => 29,
    808 => 29,
    809 => 29,
    810 => 29,
    811 => 29,
    812 => 29,
    813 => 29,
    814 => 29,
    815 => 29,
    816 => 29,
    817 => 29,
    818 => 29,
    819 => 29,
    820 => 29,
    821 => 30,
    822 => 30,
    823 => 30,
    824 => 30,
    825 => 30,
    826 => 30,
    827 => 30,
    828 => 30,
    829 => 30,
    830 => 30,
    831 => 30,
    832 => 30,
    833 => 30,
    834 => 30,
    835 => 30,
    836 => 30,
    837 => 30,
    838 => 30,
    839 => 30,
    840 => 30,
    841 => 30,
    842 => 30,
    843 => 30,
    844 => 30,
    845 => 30,
    846 => 30,
    847 => 30,
    848 => 30,
    849 => 30,
    850 => 30,
    851 => 30,
    852 => 30,
    853 => 30,
    854 => 30,
    855 => 30,
    856 => 30,
    857 => 30,
    858 => 30,
    859 => 30,
    860 => 30,
    861 => 30,
    862 => 30,
    863 => 30,
    864 => 30,
    865 => 30,
    866 => 30,
    867 => 30,
    868 => 30,
    869 => 30,
    870 => 30,
    871 => 30,
    872 => 30,
    873 => 30,
    874 => 30,
    875 => 30,
    876 => 30,
    877 => 30,
    878 => 30,
    879 => 30,
    880 => 30,
    881 => 30,
    882 => 30,
    883 => 30,
    884 => 30,
    885 => 30,
    886 => 30,
    887 => 30,
    888 => 30,
    889 => 30,
    890 => 30,
    891 => 30,
    892 => 30,
    893 => 30,
    894 => 30,
    895 => 30,
    896 => 30,
    897 => 30,
    898 => 30,
    899 => 30,
    900 => 30,
    901 => 30,
    902 => 30,
    903 => 30,
    904 => 30,
    905 => 30,
    906 => 30,
    907 => 31,
    908 => 31,
    909 => 31,
    910 => 31,
    911 => 31,
    912 => 31,
    913 => 31,
    914 => 31,
    915 => 31,
    916 => 31,
    917 => 31,
    918 => 31,
    919 => 31,
    920 => 31,
    921 => 31,
    922 => 31,
    923 => 31,
    924 => 31,
    925 => 31,
    926 => 31,
    927 => 31,
    928 => 31,
    929 => 31,
    930 => 31,
    931 => 31,
    932 => 31,
    933 => 31,
    934 => 31,
    935 => 31,
    936 => 31,
    937 => 31,
    938 => 31,
    939 => 31,
    940 => 31,
    941 => 31,
    942 => 31,
    943 => 31,
    944 => 31,
    945 => 31,
    946 => 31,
    947 => 31,
    948 => 31,
    949 => 31,
    950 => 31,
    951 => 31,
    952 => 31,
    953 => 31,
    954 => 31,
    955 => 31,
    956 => 31,
    957 => 31,
    958 => 31,
    959 => 31,
    960 => 31,
    961 => 31,
    962 => 31,
    963 => 31,
    964 => 31,
    965 => 31,
    966 => 31,
    967 => 31,
    968 => 31,
    969 => 31,
    970 => 31,
    971 => 31,
    972 => 31,
    973 => 31,
    974 => 31,
    975 => 31,
    976 => 31,
    977 => 31,
    978 => 31,
    979 => 31,
    980 => 31,
    981 => 31,
    982 => 31,
    983 => 31,
    984 => 31,
    985 => 31,
    986 => 31,
    987 => 31,
    988 => 31,
    989 => 31,
    990 => 31,
    991 => 31,
    992 => 31,
    993 => 31,
    994 => 31,
    995 => 31,
    996 => 31,
    997 => 31,
    998 => 31,
    999 => 31,
    1000 => 31,
    1001 => 31,
    1002 => 31,
    1003 => 31,
    1004 => 31,
    1005 => 31,
    1006 => 31,
    1007 => 31,
    1008 => 31,
    1009 => 31,
    1010 => 31,
    1011 => 31,
    1012 => 31,
    1013 => 31,
    1014 => 31,
    1015 => 31,
    1016 => 31,
    1017 => 31,
    1018 => 31,
    1019 => 31,
    1020 => 31,
    1021 => 31,
    1022 => 31,
    1023 => 31,
    1024 => 31,
    1025 => 31,
    1026 => 31,
    1027 => 31,
    1028 => 31,
    1029 => 31,
    1030 => 31,
    1031 => 31,
    1032 => 31,
    1033 => 31,
    1034 => 31,
    1035 => 31,
    1036 => 31,
    1037 => 31,
    1038 => 31,
    1039 => 31,
    1040 => 31,
    1041 => 31,
    1042 => 31,
    1043 => 31,
    1044 => 31,
    1045 => 31,
    1046 => 31,
    1047 => 31,
    1048 => 31,
    1049 => 31,
    1050 => 31,
    1051 => 31,
    1052 => 31,
    1053 => 31,
    1054 => 31,
    1055 => 31,
    1056 => 31,
    1057 => 31,
    1058 => 31,
    1059 => 31,
    1060 => 31,
    1061 => 31,
    1062 => 31,
    1063 => 31,
    1064 => 31,
    1065 => 31,
    1066 => 31,
    1067 => 31,
    1068 => 31,
    1069 => 31,
    1070 => 31,
    1071 => 31,
    1072 => 31,
    1073 => 31,
    1074 => 31,
    1075 => 31,
    1076 => 31,
    1077 => 31,
    1078 => 31,
    1079 => 31,
    1080 => 31,
    1081 => 31,
    1082 => 31,
    1083 => 31,
    1084 => 31,
    1085 => 31,
    1086 => 31,
    1087 => 31,
    1088 => 31,
    1089 => 31,
    1090 => 31,
    1091 => 31,
    1092 => 31,
    1093 => 31,
    1094 => 31,
    1095 => 31,
    1096 => 31,
    1097 => 31,
    1098 => 31,
    1099 => 31,
    1100 => 31,
    1101 => 31,
    1102 => 31,
    1103 => 31,
    1104 => 31,
    1105 => 31,
    1106 => 31,
    1107 => 31,
    1108 => 31,
    1109 => 31,
    1110 => 31,
    1111 => 31,
    1112 => 31,
    1113 => 31,
    1114 => 31,
    1115 => 31,
    1116 => 31,
    1117 => 31,
    1118 => 31,
    1119 => 31,
    1120 => 31,
    1121 => 31,
    1122 => 31,
    1123 => 31,
    1124 => 31,
    1125 => 31,
    1126 => 31,
    1127 => 31,
    1128 => 31,
    1129 => 31,
    1130 => 31,
    1131 => 31,
    1132 => 31,
    1133 => 31,
    1134 => 31,
    1135 => 31,
    1136 => 31,
    1137 => 31,
    1138 => 31,
    1139 => 31,
    1140 => 31,
    1141 => 31,
    1142 => 30,
    1143 => 30,
    1144 => 30,
    1145 => 30,
    1146 => 30,
    1147 => 30,
    1148 => 30,
    1149 => 30,
    1150 => 30,
    1151 => 30,
    1152 => 30,
    1153 => 30,
    1154 => 30,
    1155 => 30,
    1156 => 30,
    1157 => 30,
    1158 => 30,
    1159 => 30,
    1160 => 30,
    1161 => 30,
    1162 => 30,
    1163 => 30,
    1164 => 30,
    1165 => 30,
    1166 => 30,
    1167 => 30,
    1168 => 30,
    1169 => 30,
    1170 => 30,
    1171 => 30,
    1172 => 30,
    1173 => 30,
    1174 => 30,
    1175 => 30,
    1176 => 30,
    1177 => 30,
    1178 => 30,
    1179 => 30,
    1180 => 30,
    1181 => 30,
    1182 => 30,
    1183 => 30,
    1184 => 30,
    1185 => 30,
    1186 => 30,
    1187 => 30,
    1188 => 30,
    1189 => 30,
    1190 => 30,
    1191 => 30,
    1192 => 30,
    1193 => 30,
    1194 => 30,
    1195 => 30,
    1196 => 30,
    1197 => 30,
    1198 => 30,
    1199 => 30,
    1200 => 30,
    1201 => 30,
    1202 => 30,
    1203 => 30,
    1204 => 30,
    1205 => 30,
    1206 => 30,
    1207 => 30,
    1208 => 30,
    1209 => 30,
    1210 => 30,
    1211 => 30,
    1212 => 30,
    1213 => 30,
    1214 => 30,
    1215 => 30,
    1216 => 30,
    1217 => 30,
    1218 => 30,
    1219 => 30,
    1220 => 30,
    1221 => 30,
    1222 => 30,
    1223 => 30,
    1224 => 30,
    1225 => 30,
    1226 => 30,
    1227 => 30,
    1228 => 29,
    1229 => 29,
    1230 => 29,
    1231 => 29,
    1232 => 29,
    1233 => 29,
    1234 => 29,
    1235 => 29,
    1236 => 29,
    1237 => 29,
    1238 => 29,
    1239 => 29,
    1240 => 29,
    1241 => 29,
    1242 => 29,
    1243 => 29,
    1244 => 29,
    1245 => 29,
    1246 => 29,
    1247 => 29,
    1248 => 29,
    1249 => 29,
    1250 => 29,
    1251 => 29,
    1252 => 29,
    1253 => 29,
    1254 => 29,
    1255 => 29,
    1256 => 29,
    1257 => 29,
    1258 => 29,
    1259 => 29,
    1260 => 29,
    1261 => 29,
    1262 => 29,
    1263 => 29,
    1264 => 29,
    1265 => 29,
    1266 => 29,
    1267 => 29,
    1268 => 29,
    1269 => 29,
    1270 => 29,
    1271 => 29,
    1272 => 29,
    1273 => 29,
    1274 => 29,
    1275 => 29,
    1276 => 29,
    1277 => 29,
    1278 => 29,
    1279 => 29,
    1280 => 29,
    1281 => 29,
    1282 => 29,
    1283 => 29,
    1284 => 29,
    1285 => 29,
    1286 => 29,
    1287 => 29,
    1288 => 28,
    1289 => 28,
    1290 => 28,
    1291 => 28,
    1292 => 28,
    1293 => 28,
    1294 => 28,
    1295 => 28,
    1296 => 28,
    1297 => 28,
    1298 => 28,
    1299 => 28,
    1300 => 28,
    1301 => 28,
    1302 => 28,
    1303 => 28,
    1304 => 28,
    1305 => 28,
    1306 => 28,
    1307 => 28,
    1308 => 28,
    1309 => 28,
    1310 => 28,
    1311 => 28,
    1312 => 28,
    1313 => 28,
    1314 => 28,
    1315 => 28,
    1316 => 28,
    1317 => 28,
    1318 => 28,
    1319 => 28,
    1320 => 28,
    1321 => 28,
    1322 => 28,
    1323 => 28,
    1324 => 28,
    1325 => 28,
    1326 => 28,
    1327 => 28,
    1328 => 28,
    1329 => 28,
    1330 => 28,
    1331 => 28,
    1332 => 28,
    1333 => 28,
    1334 => 28,
    1335 => 28,
    1336 => 28,
    1337 => 27,
    1338 => 27,
    1339 => 27,
    1340 => 27,
    1341 => 27,
    1342 => 27,
    1343 => 27,
    1344 => 27,
    1345 => 27,
    1346 => 27,
    1347 => 27,
    1348 => 27,
    1349 => 27,
    1350 => 27,
    1351 => 27,
    1352 => 27,
    1353 => 27,
    1354 => 27,
    1355 => 27,
    1356 => 27,
    1357 => 27,
    1358 => 27,
    1359 => 27,
    1360 => 27,
    1361 => 27,
    1362 => 27,
    1363 => 27,
    1364 => 27,
    1365 => 27,
    1366 => 27,
    1367 => 27,
    1368 => 27,
    1369 => 27,
    1370 => 27,
    1371 => 27,
    1372 => 27,
    1373 => 27,
    1374 => 27,
    1375 => 27,
    1376 => 27,
    1377 => 27,
    1378 => 27,
    1379 => 27,
    1380 => 26,
    1381 => 26,
    1382 => 26,
    1383 => 26,
    1384 => 26,
    1385 => 26,
    1386 => 26,
    1387 => 26,
    1388 => 26,
    1389 => 26,
    1390 => 26,
    1391 => 26,
    1392 => 26,
    1393 => 26,
    1394 => 26,
    1395 => 26,
    1396 => 26,
    1397 => 26,
    1398 => 26,
    1399 => 26,
    1400 => 26,
    1401 => 26,
    1402 => 26,
    1403 => 26,
    1404 => 26,
    1405 => 26,
    1406 => 26,
    1407 => 26,
    1408 => 26,
    1409 => 26,
    1410 => 26,
    1411 => 26,
    1412 => 26,
    1413 => 26,
    1414 => 26,
    1415 => 26,
    1416 => 26,
    1417 => 26,
    1418 => 26,
    1419 => 25,
    1420 => 25,
    1421 => 25,
    1422 => 25,
    1423 => 25,
    1424 => 25,
    1425 => 25,
    1426 => 25,
    1427 => 25,
    1428 => 25,
    1429 => 25,
    1430 => 25,
    1431 => 25,
    1432 => 25,
    1433 => 25,
    1434 => 25,
    1435 => 25,
    1436 => 25,
    1437 => 25,
    1438 => 25,
    1439 => 25,
    1440 => 25,
    1441 => 25,
    1442 => 25,
    1443 => 25,
    1444 => 25,
    1445 => 25,
    1446 => 25,
    1447 => 25,
    1448 => 25,
    1449 => 25,
    1450 => 25,
    1451 => 25,
    1452 => 25,
    1453 => 25,
    1454 => 24,
    1455 => 24,
    1456 => 24,
    1457 => 24,
    1458 => 24,
    1459 => 24,
    1460 => 24,
    1461 => 24,
    1462 => 24,
    1463 => 24,
    1464 => 24,
    1465 => 24,
    1466 => 24,
    1467 => 24,
    1468 => 24,
    1469 => 24,
    1470 => 24,
    1471 => 24,
    1472 => 24,
    1473 => 24,
    1474 => 24,
    1475 => 24,
    1476 => 24,
    1477 => 24,
    1478 => 24,
    1479 => 24,
    1480 => 24,
    1481 => 24,
    1482 => 24,
    1483 => 24,
    1484 => 24,
    1485 => 24,
    1486 => 24,
    1487 => 24,
    1488 => 23,
    1489 => 23,
    1490 => 23,
    1491 => 23,
    1492 => 23,
    1493 => 23,
    1494 => 23,
    1495 => 23,
    1496 => 23,
    1497 => 23,
    1498 => 23,
    1499 => 23,
    1500 => 23,
    1501 => 23,
    1502 => 23,
    1503 => 23,
    1504 => 23,
    1505 => 23,
    1506 => 23,
    1507 => 23,
    1508 => 23,
    1509 => 23,
    1510 => 23,
    1511 => 23,
    1512 => 23,
    1513 => 23,
    1514 => 23,
    1515 => 23,
    1516 => 23,
    1517 => 23,
    1518 => 23,
    1519 => 22,
    1520 => 22,
    1521 => 22,
    1522 => 22,
    1523 => 22,
    1524 => 22,
    1525 => 22,
    1526 => 22,
    1527 => 22,
    1528 => 22,
    1529 => 22,
    1530 => 22,
    1531 => 22,
    1532 => 22,
    1533 => 22,
    1534 => 22,
    1535 => 22,
    1536 => 22,
    1537 => 22,
    1538 => 22,
    1539 => 22,
    1540 => 22,
    1541 => 22,
    1542 => 22,
    1543 => 22,
    1544 => 22,
    1545 => 22,
    1546 => 22,
    1547 => 22,
    1548 => 22,
    1549 => 21,
    1550 => 21,
    1551 => 21,
    1552 => 21,
    1553 => 21,
    1554 => 21,
    1555 => 21,
    1556 => 21,
    1557 => 21,
    1558 => 21,
    1559 => 21,
    1560 => 21,
    1561 => 21,
    1562 => 21,
    1563 => 21,
    1564 => 21,
    1565 => 21,
    1566 => 21,
    1567 => 21,
    1568 => 21,
    1569 => 21,
    1570 => 21,
    1571 => 21,
    1572 => 21,
    1573 => 21,
    1574 => 21,
    1575 => 21,
    1576 => 21,
    1577 => 20,
    1578 => 20,
    1579 => 20,
    1580 => 20,
    1581 => 20,
    1582 => 20,
    1583 => 20,
    1584 => 20,
    1585 => 20,
    1586 => 20,
    1587 => 20,
    1588 => 20,
    1589 => 20,
    1590 => 20,
    1591 => 20,
    1592 => 20,
    1593 => 20,
    1594 => 20,
    1595 => 20,
    1596 => 20,
    1597 => 20,
    1598 => 20,
    1599 => 20,
    1600 => 20,
    1601 => 20,
    1602 => 20,
    1603 => 20,
    1604 => 20,
    1605 => 19,
    1606 => 19,
    1607 => 19,
    1608 => 19,
    1609 => 19,
    1610 => 19,
    1611 => 19,
    1612 => 19,
    1613 => 19,
    1614 => 19,
    1615 => 19,
    1616 => 19,
    1617 => 19,
    1618 => 19,
    1619 => 19,
    1620 => 19,
    1621 => 19,
    1622 => 19,
    1623 => 19,
    1624 => 19,
    1625 => 19,
    1626 => 19,
    1627 => 19,
    1628 => 19,
    1629 => 19,
    1630 => 19,
    1631 => 19,
    1632 => 18,
    1633 => 18,
    1634 => 18,
    1635 => 18,
    1636 => 18,
    1637 => 18,
    1638 => 18,
    1639 => 18,
    1640 => 18,
    1641 => 18,
    1642 => 18,
    1643 => 18,
    1644 => 18,
    1645 => 18,
    1646 => 18,
    1647 => 18,
    1648 => 18,
    1649 => 18,
    1650 => 18,
    1651 => 18,
    1652 => 18,
    1653 => 18,
    1654 => 18,
    1655 => 18,
    1656 => 18,
    1657 => 17,
    1658 => 17,
    1659 => 17,
    1660 => 17,
    1661 => 17,
    1662 => 17,
    1663 => 17,
    1664 => 17,
    1665 => 17,
    1666 => 17,
    1667 => 17,
    1668 => 17,
    1669 => 17,
    1670 => 17,
    1671 => 17,
    1672 => 17,
    1673 => 17,
    1674 => 17,
    1675 => 17,
    1676 => 17,
    1677 => 17,
    1678 => 17,
    1679 => 17,
    1680 => 17,
    1681 => 17,
    1682 => 17,
    1683 => 16,
    1684 => 16,
    1685 => 16,
    1686 => 16,
    1687 => 16,
    1688 => 16,
    1689 => 16,
    1690 => 16,
    1691 => 16,
    1692 => 16,
    1693 => 16,
    1694 => 16,
    1695 => 16,
    1696 => 16,
    1697 => 16,
    1698 => 16,
    1699 => 16,
    1700 => 16,
    1701 => 16,
    1702 => 16,
    1703 => 16,
    1704 => 16,
    1705 => 16,
    1706 => 16,
    1707 => 15,
    1708 => 15,
    1709 => 15,
    1710 => 15,
    1711 => 15,
    1712 => 15,
    1713 => 15,
    1714 => 15,
    1715 => 15,
    1716 => 15,
    1717 => 15,
    1718 => 15,
    1719 => 15,
    1720 => 15,
    1721 => 15,
    1722 => 15,
    1723 => 15,
    1724 => 15,
    1725 => 15,
    1726 => 15,
    1727 => 15,
    1728 => 15,
    1729 => 15,
    1730 => 15,
    1731 => 14,
    1732 => 14,
    1733 => 14,
    1734 => 14,
    1735 => 14,
    1736 => 14,
    1737 => 14,
    1738 => 14,
    1739 => 14,
    1740 => 14,
    1741 => 14,
    1742 => 14,
    1743 => 14,
    1744 => 14,
    1745 => 14,
    1746 => 14,
    1747 => 14,
    1748 => 14,
    1749 => 14,
    1750 => 14,
    1751 => 14,
    1752 => 14,
    1753 => 14,
    1754 => 14,
    1755 => 13,
    1756 => 13,
    1757 => 13,
    1758 => 13,
    1759 => 13,
    1760 => 13,
    1761 => 13,
    1762 => 13,
    1763 => 13,
    1764 => 13,
    1765 => 13,
    1766 => 13,
    1767 => 13,
    1768 => 13,
    1769 => 13,
    1770 => 13,
    1771 => 13,
    1772 => 13,
    1773 => 13,
    1774 => 13,
    1775 => 13,
    1776 => 13,
    1777 => 13,
    1778 => 12,
    1779 => 12,
    1780 => 12,
    1781 => 12,
    1782 => 12,
    1783 => 12,
    1784 => 12,
    1785 => 12,
    1786 => 12,
    1787 => 12,
    1788 => 12,
    1789 => 12,
    1790 => 12,
    1791 => 12,
    1792 => 12,
    1793 => 12,
    1794 => 12,
    1795 => 12,
    1796 => 12,
    1797 => 12,
    1798 => 12,
    1799 => 12,
    1800 => 12,
    1801 => 11,
    1802 => 11,
    1803 => 11,
    1804 => 11,
    1805 => 11,
    1806 => 11,
    1807 => 11,
    1808 => 11,
    1809 => 11,
    1810 => 11,
    1811 => 11,
    1812 => 11,
    1813 => 11,
    1814 => 11,
    1815 => 11,
    1816 => 11,
    1817 => 11,
    1818 => 11,
    1819 => 11,
    1820 => 11,
    1821 => 11,
    1822 => 11,
    1823 => 10,
    1824 => 10,
    1825 => 10,
    1826 => 10,
    1827 => 10,
    1828 => 10,
    1829 => 10,
    1830 => 10,
    1831 => 10,
    1832 => 10,
    1833 => 10,
    1834 => 10,
    1835 => 10,
    1836 => 10,
    1837 => 10,
    1838 => 10,
    1839 => 10,
    1840 => 10,
    1841 => 10,
    1842 => 10,
    1843 => 10,
    1844 => 10,
    1845 => 9,
    1846 => 9,
    1847 => 9,
    1848 => 9,
    1849 => 9,
    1850 => 9,
    1851 => 9,
    1852 => 9,
    1853 => 9,
    1854 => 9,
    1855 => 9,
    1856 => 9,
    1857 => 9,
    1858 => 9,
    1859 => 9,
    1860 => 9,
    1861 => 9,
    1862 => 9,
    1863 => 9,
    1864 => 9,
    1865 => 9,
    1866 => 9,
    1867 => 8,
    1868 => 8,
    1869 => 8,
    1870 => 8,
    1871 => 8,
    1872 => 8,
    1873 => 8,
    1874 => 8,
    1875 => 8,
    1876 => 8,
    1877 => 8,
    1878 => 8,
    1879 => 8,
    1880 => 8,
    1881 => 8,
    1882 => 8,
    1883 => 8,
    1884 => 8,
    1885 => 8,
    1886 => 8,
    1887 => 8,
    1888 => 8,
    1889 => 7,
    1890 => 7,
    1891 => 7,
    1892 => 7,
    1893 => 7,
    1894 => 7,
    1895 => 7,
    1896 => 7,
    1897 => 7,
    1898 => 7,
    1899 => 7,
    1900 => 7,
    1901 => 7,
    1902 => 7,
    1903 => 7,
    1904 => 7,
    1905 => 7,
    1906 => 7,
    1907 => 7,
    1908 => 7,
    1909 => 7,
    1910 => 7,
    1911 => 6,
    1912 => 6,
    1913 => 6,
    1914 => 6,
    1915 => 6,
    1916 => 6,
    1917 => 6,
    1918 => 6,
    1919 => 6,
    1920 => 6,
    1921 => 6,
    1922 => 6,
    1923 => 6,
    1924 => 6,
    1925 => 6,
    1926 => 6,
    1927 => 6,
    1928 => 6,
    1929 => 6,
    1930 => 6,
    1931 => 6,
    1932 => 5,
    1933 => 5,
    1934 => 5,
    1935 => 5,
    1936 => 5,
    1937 => 5,
    1938 => 5,
    1939 => 5,
    1940 => 5,
    1941 => 5,
    1942 => 5,
    1943 => 5,
    1944 => 5,
    1945 => 5,
    1946 => 5,
    1947 => 5,
    1948 => 5,
    1949 => 5,
    1950 => 5,
    1951 => 5,
    1952 => 5,
    1953 => 5,
    1954 => 4,
    1955 => 4,
    1956 => 4,
    1957 => 4,
    1958 => 4,
    1959 => 4,
    1960 => 4,
    1961 => 4,
    1962 => 4,
    1963 => 4,
    1964 => 4,
    1965 => 4,
    1966 => 4,
    1967 => 4,
    1968 => 4,
    1969 => 4,
    1970 => 4,
    1971 => 4,
    1972 => 4,
    1973 => 4,
    1974 => 4,
    1975 => 3,
    1976 => 3,
    1977 => 3,
    1978 => 3,
    1979 => 3,
    1980 => 3,
    1981 => 3,
    1982 => 3,
    1983 => 3,
    1984 => 3,
    1985 => 3,
    1986 => 3,
    1987 => 3,
    1988 => 3,
    1989 => 3,
    1990 => 3,
    1991 => 3,
    1992 => 3,
    1993 => 3,
    1994 => 3,
    1995 => 3,
    1996 => 2,
    1997 => 2,
    1998 => 2,
    1999 => 2,
    2000 => 2,
    2001 => 2,
    2002 => 2,
    2003 => 2,
    2004 => 2,
    2005 => 2,
    2006 => 2,
    2007 => 2,
    2008 => 2,
    2009 => 2,
    2010 => 2,
    2011 => 2,
    2012 => 2,
    2013 => 2,
    2014 => 2,
    2015 => 2,
    2016 => 2,
    2017 => 1,
    2018 => 1,
    2019 => 1,
    2020 => 1,
    2021 => 1,
    2022 => 1,
    2023 => 1,
    2024 => 1,
    2025 => 1,
    2026 => 1,
    2027 => 1,
    2028 => 1,
    2029 => 1,
    2030 => 1,
    2031 => 1,
    2032 => 1,
    2033 => 1,
    2034 => 1,
    2035 => 1,
    2036 => 1,
    2037 => 1,
    2038 => 0,
    2039 => 0,
    2040 => 0,
    2041 => 0,
    2042 => 0,
    2043 => 0,
    2044 => 0,
    2045 => 0,
    2046 => 0,
    2047 => 0,
    2048 => 0,
    2049 => 0,
    2050 => 0,
    2051 => 0,
    2052 => 0,
    2053 => 0,
    2054 => 0,
    2055 => 0,
    2056 => 0,
    2057 => 0,
    2058 => 0,
    2059 => -1,
    2060 => -1,
    2061 => -1,
    2062 => -1,
    2063 => -1,
    2064 => -1,
    2065 => -1,
    2066 => -1,
    2067 => -1,
    2068 => -1,
    2069 => -1,
    2070 => -1,
    2071 => -1,
    2072 => -1,
    2073 => -1,
    2074 => -1,
    2075 => -1,
    2076 => -1,
    2077 => -1,
    2078 => -1,
    2079 => -1,
    2080 => -2,
    2081 => -2,
    2082 => -2,
    2083 => -2,
    2084 => -2,
    2085 => -2,
    2086 => -2,
    2087 => -2,
    2088 => -2,
    2089 => -2,
    2090 => -2,
    2091 => -2,
    2092 => -2,
    2093 => -2,
    2094 => -2,
    2095 => -2,
    2096 => -2,
    2097 => -2,
    2098 => -2,
    2099 => -2,
    2100 => -2,
    2101 => -3,
    2102 => -3,
    2103 => -3,
    2104 => -3,
    2105 => -3,
    2106 => -3,
    2107 => -3,
    2108 => -3,
    2109 => -3,
    2110 => -3,
    2111 => -3,
    2112 => -3,
    2113 => -3,
    2114 => -3,
    2115 => -3,
    2116 => -3,
    2117 => -3,
    2118 => -3,
    2119 => -3,
    2120 => -3,
    2121 => -3,
    2122 => -4,
    2123 => -4,
    2124 => -4,
    2125 => -4,
    2126 => -4,
    2127 => -4,
    2128 => -4,
    2129 => -4,
    2130 => -4,
    2131 => -4,
    2132 => -4,
    2133 => -4,
    2134 => -4,
    2135 => -4,
    2136 => -4,
    2137 => -4,
    2138 => -4,
    2139 => -4,
    2140 => -4,
    2141 => -4,
    2142 => -4,
    2143 => -5,
    2144 => -5,
    2145 => -5,
    2146 => -5,
    2147 => -5,
    2148 => -5,
    2149 => -5,
    2150 => -5,
    2151 => -5,
    2152 => -5,
    2153 => -5,
    2154 => -5,
    2155 => -5,
    2156 => -5,
    2157 => -5,
    2158 => -5,
    2159 => -5,
    2160 => -5,
    2161 => -5,
    2162 => -5,
    2163 => -5,
    2164 => -5,
    2165 => -6,
    2166 => -6,
    2167 => -6,
    2168 => -6,
    2169 => -6,
    2170 => -6,
    2171 => -6,
    2172 => -6,
    2173 => -6,
    2174 => -6,
    2175 => -6,
    2176 => -6,
    2177 => -6,
    2178 => -6,
    2179 => -6,
    2180 => -6,
    2181 => -6,
    2182 => -6,
    2183 => -6,
    2184 => -6,
    2185 => -6,
    2186 => -7,
    2187 => -7,
    2188 => -7,
    2189 => -7,
    2190 => -7,
    2191 => -7,
    2192 => -7,
    2193 => -7,
    2194 => -7,
    2195 => -7,
    2196 => -7,
    2197 => -7,
    2198 => -7,
    2199 => -7,
    2200 => -7,
    2201 => -7,
    2202 => -7,
    2203 => -7,
    2204 => -7,
    2205 => -7,
    2206 => -7,
    2207 => -7,
    2208 => -8,
    2209 => -8,
    2210 => -8,
    2211 => -8,
    2212 => -8,
    2213 => -8,
    2214 => -8,
    2215 => -8,
    2216 => -8,
    2217 => -8,
    2218 => -8,
    2219 => -8,
    2220 => -8,
    2221 => -8,
    2222 => -8,
    2223 => -8,
    2224 => -8,
    2225 => -8,
    2226 => -8,
    2227 => -8,
    2228 => -8,
    2229 => -8,
    2230 => -9,
    2231 => -9,
    2232 => -9,
    2233 => -9,
    2234 => -9,
    2235 => -9,
    2236 => -9,
    2237 => -9,
    2238 => -9,
    2239 => -9,
    2240 => -9,
    2241 => -9,
    2242 => -9,
    2243 => -9,
    2244 => -9,
    2245 => -9,
    2246 => -9,
    2247 => -9,
    2248 => -9,
    2249 => -9,
    2250 => -9,
    2251 => -9,
    2252 => -10,
    2253 => -10,
    2254 => -10,
    2255 => -10,
    2256 => -10,
    2257 => -10,
    2258 => -10,
    2259 => -10,
    2260 => -10,
    2261 => -10,
    2262 => -10,
    2263 => -10,
    2264 => -10,
    2265 => -10,
    2266 => -10,
    2267 => -10,
    2268 => -10,
    2269 => -10,
    2270 => -10,
    2271 => -10,
    2272 => -10,
    2273 => -10,
    2274 => -11,
    2275 => -11,
    2276 => -11,
    2277 => -11,
    2278 => -11,
    2279 => -11,
    2280 => -11,
    2281 => -11,
    2282 => -11,
    2283 => -11,
    2284 => -11,
    2285 => -11,
    2286 => -11,
    2287 => -11,
    2288 => -11,
    2289 => -11,
    2290 => -11,
    2291 => -11,
    2292 => -11,
    2293 => -11,
    2294 => -11,
    2295 => -11,
    2296 => -12,
    2297 => -12,
    2298 => -12,
    2299 => -12,
    2300 => -12,
    2301 => -12,
    2302 => -12,
    2303 => -12,
    2304 => -12,
    2305 => -12,
    2306 => -12,
    2307 => -12,
    2308 => -12,
    2309 => -12,
    2310 => -12,
    2311 => -12,
    2312 => -12,
    2313 => -12,
    2314 => -12,
    2315 => -12,
    2316 => -12,
    2317 => -12,
    2318 => -12,
    2319 => -13,
    2320 => -13,
    2321 => -13,
    2322 => -13,
    2323 => -13,
    2324 => -13,
    2325 => -13,
    2326 => -13,
    2327 => -13,
    2328 => -13,
    2329 => -13,
    2330 => -13,
    2331 => -13,
    2332 => -13,
    2333 => -13,
    2334 => -13,
    2335 => -13,
    2336 => -13,
    2337 => -13,
    2338 => -13,
    2339 => -13,
    2340 => -13,
    2341 => -13,
    2342 => -14,
    2343 => -14,
    2344 => -14,
    2345 => -14,
    2346 => -14,
    2347 => -14,
    2348 => -14,
    2349 => -14,
    2350 => -14,
    2351 => -14,
    2352 => -14,
    2353 => -14,
    2354 => -14,
    2355 => -14,
    2356 => -14,
    2357 => -14,
    2358 => -14,
    2359 => -14,
    2360 => -14,
    2361 => -14,
    2362 => -14,
    2363 => -14,
    2364 => -14,
    2365 => -14,
    2366 => -15,
    2367 => -15,
    2368 => -15,
    2369 => -15,
    2370 => -15,
    2371 => -15,
    2372 => -15,
    2373 => -15,
    2374 => -15,
    2375 => -15,
    2376 => -15,
    2377 => -15,
    2378 => -15,
    2379 => -15,
    2380 => -15,
    2381 => -15,
    2382 => -15,
    2383 => -15,
    2384 => -15,
    2385 => -15,
    2386 => -15,
    2387 => -15,
    2388 => -15,
    2389 => -15,
    2390 => -16,
    2391 => -16,
    2392 => -16,
    2393 => -16,
    2394 => -16,
    2395 => -16,
    2396 => -16,
    2397 => -16,
    2398 => -16,
    2399 => -16,
    2400 => -16,
    2401 => -16,
    2402 => -16,
    2403 => -16,
    2404 => -16,
    2405 => -16,
    2406 => -16,
    2407 => -16,
    2408 => -16,
    2409 => -16,
    2410 => -16,
    2411 => -16,
    2412 => -16,
    2413 => -16,
    2414 => -17,
    2415 => -17,
    2416 => -17,
    2417 => -17,
    2418 => -17,
    2419 => -17,
    2420 => -17,
    2421 => -17,
    2422 => -17,
    2423 => -17,
    2424 => -17,
    2425 => -17,
    2426 => -17,
    2427 => -17,
    2428 => -17,
    2429 => -17,
    2430 => -17,
    2431 => -17,
    2432 => -17,
    2433 => -17,
    2434 => -17,
    2435 => -17,
    2436 => -17,
    2437 => -17,
    2438 => -17,
    2439 => -17,
    2440 => -18,
    2441 => -18,
    2442 => -18,
    2443 => -18,
    2444 => -18,
    2445 => -18,
    2446 => -18,
    2447 => -18,
    2448 => -18,
    2449 => -18,
    2450 => -18,
    2451 => -18,
    2452 => -18,
    2453 => -18,
    2454 => -18,
    2455 => -18,
    2456 => -18,
    2457 => -18,
    2458 => -18,
    2459 => -18,
    2460 => -18,
    2461 => -18,
    2462 => -18,
    2463 => -18,
    2464 => -18,
    2465 => -19,
    2466 => -19,
    2467 => -19,
    2468 => -19,
    2469 => -19,
    2470 => -19,
    2471 => -19,
    2472 => -19,
    2473 => -19,
    2474 => -19,
    2475 => -19,
    2476 => -19,
    2477 => -19,
    2478 => -19,
    2479 => -19,
    2480 => -19,
    2481 => -19,
    2482 => -19,
    2483 => -19,
    2484 => -19,
    2485 => -19,
    2486 => -19,
    2487 => -19,
    2488 => -19,
    2489 => -19,
    2490 => -19,
    2491 => -19,
    2492 => -20,
    2493 => -20,
    2494 => -20,
    2495 => -20,
    2496 => -20,
    2497 => -20,
    2498 => -20,
    2499 => -20,
    2500 => -20,
    2501 => -20,
    2502 => -20,
    2503 => -20,
    2504 => -20,
    2505 => -20,
    2506 => -20,
    2507 => -20,
    2508 => -20,
    2509 => -20,
    2510 => -20,
    2511 => -20,
    2512 => -20,
    2513 => -20,
    2514 => -20,
    2515 => -20,
    2516 => -20,
    2517 => -20,
    2518 => -20,
    2519 => -20,
    2520 => -21,
    2521 => -21,
    2522 => -21,
    2523 => -21,
    2524 => -21,
    2525 => -21,
    2526 => -21,
    2527 => -21,
    2528 => -21,
    2529 => -21,
    2530 => -21,
    2531 => -21,
    2532 => -21,
    2533 => -21,
    2534 => -21,
    2535 => -21,
    2536 => -21,
    2537 => -21,
    2538 => -21,
    2539 => -21,
    2540 => -21,
    2541 => -21,
    2542 => -21,
    2543 => -21,
    2544 => -21,
    2545 => -21,
    2546 => -21,
    2547 => -21,
    2548 => -22,
    2549 => -22,
    2550 => -22,
    2551 => -22,
    2552 => -22,
    2553 => -22,
    2554 => -22,
    2555 => -22,
    2556 => -22,
    2557 => -22,
    2558 => -22,
    2559 => -22,
    2560 => -22,
    2561 => -22,
    2562 => -22,
    2563 => -22,
    2564 => -22,
    2565 => -22,
    2566 => -22,
    2567 => -22,
    2568 => -22,
    2569 => -22,
    2570 => -22,
    2571 => -22,
    2572 => -22,
    2573 => -22,
    2574 => -22,
    2575 => -22,
    2576 => -22,
    2577 => -22,
    2578 => -23,
    2579 => -23,
    2580 => -23,
    2581 => -23,
    2582 => -23,
    2583 => -23,
    2584 => -23,
    2585 => -23,
    2586 => -23,
    2587 => -23,
    2588 => -23,
    2589 => -23,
    2590 => -23,
    2591 => -23,
    2592 => -23,
    2593 => -23,
    2594 => -23,
    2595 => -23,
    2596 => -23,
    2597 => -23,
    2598 => -23,
    2599 => -23,
    2600 => -23,
    2601 => -23,
    2602 => -23,
    2603 => -23,
    2604 => -23,
    2605 => -23,
    2606 => -23,
    2607 => -23,
    2608 => -23,
    2609 => -24,
    2610 => -24,
    2611 => -24,
    2612 => -24,
    2613 => -24,
    2614 => -24,
    2615 => -24,
    2616 => -24,
    2617 => -24,
    2618 => -24,
    2619 => -24,
    2620 => -24,
    2621 => -24,
    2622 => -24,
    2623 => -24,
    2624 => -24,
    2625 => -24,
    2626 => -24,
    2627 => -24,
    2628 => -24,
    2629 => -24,
    2630 => -24,
    2631 => -24,
    2632 => -24,
    2633 => -24,
    2634 => -24,
    2635 => -24,
    2636 => -24,
    2637 => -24,
    2638 => -24,
    2639 => -24,
    2640 => -24,
    2641 => -24,
    2642 => -24,
    2643 => -25,
    2644 => -25,
    2645 => -25,
    2646 => -25,
    2647 => -25,
    2648 => -25,
    2649 => -25,
    2650 => -25,
    2651 => -25,
    2652 => -25,
    2653 => -25,
    2654 => -25,
    2655 => -25,
    2656 => -25,
    2657 => -25,
    2658 => -25,
    2659 => -25,
    2660 => -25,
    2661 => -25,
    2662 => -25,
    2663 => -25,
    2664 => -25,
    2665 => -25,
    2666 => -25,
    2667 => -25,
    2668 => -25,
    2669 => -25,
    2670 => -25,
    2671 => -25,
    2672 => -25,
    2673 => -25,
    2674 => -25,
    2675 => -25,
    2676 => -25,
    2677 => -25,
    2678 => -26,
    2679 => -26,
    2680 => -26,
    2681 => -26,
    2682 => -26,
    2683 => -26,
    2684 => -26,
    2685 => -26,
    2686 => -26,
    2687 => -26,
    2688 => -26,
    2689 => -26,
    2690 => -26,
    2691 => -26,
    2692 => -26,
    2693 => -26,
    2694 => -26,
    2695 => -26,
    2696 => -26,
    2697 => -26,
    2698 => -26,
    2699 => -26,
    2700 => -26,
    2701 => -26,
    2702 => -26,
    2703 => -26,
    2704 => -26,
    2705 => -26,
    2706 => -26,
    2707 => -26,
    2708 => -26,
    2709 => -26,
    2710 => -26,
    2711 => -26,
    2712 => -26,
    2713 => -26,
    2714 => -26,
    2715 => -26,
    2716 => -26,
    2717 => -27,
    2718 => -27,
    2719 => -27,
    2720 => -27,
    2721 => -27,
    2722 => -27,
    2723 => -27,
    2724 => -27,
    2725 => -27,
    2726 => -27,
    2727 => -27,
    2728 => -27,
    2729 => -27,
    2730 => -27,
    2731 => -27,
    2732 => -27,
    2733 => -27,
    2734 => -27,
    2735 => -27,
    2736 => -27,
    2737 => -27,
    2738 => -27,
    2739 => -27,
    2740 => -27,
    2741 => -27,
    2742 => -27,
    2743 => -27,
    2744 => -27,
    2745 => -27,
    2746 => -27,
    2747 => -27,
    2748 => -27,
    2749 => -27,
    2750 => -27,
    2751 => -27,
    2752 => -27,
    2753 => -27,
    2754 => -27,
    2755 => -27,
    2756 => -27,
    2757 => -27,
    2758 => -27,
    2759 => -27,
    2760 => -28,
    2761 => -28,
    2762 => -28,
    2763 => -28,
    2764 => -28,
    2765 => -28,
    2766 => -28,
    2767 => -28,
    2768 => -28,
    2769 => -28,
    2770 => -28,
    2771 => -28,
    2772 => -28,
    2773 => -28,
    2774 => -28,
    2775 => -28,
    2776 => -28,
    2777 => -28,
    2778 => -28,
    2779 => -28,
    2780 => -28,
    2781 => -28,
    2782 => -28,
    2783 => -28,
    2784 => -28,
    2785 => -28,
    2786 => -28,
    2787 => -28,
    2788 => -28,
    2789 => -28,
    2790 => -28,
    2791 => -28,
    2792 => -28,
    2793 => -28,
    2794 => -28,
    2795 => -28,
    2796 => -28,
    2797 => -28,
    2798 => -28,
    2799 => -28,
    2800 => -28,
    2801 => -28,
    2802 => -28,
    2803 => -28,
    2804 => -28,
    2805 => -28,
    2806 => -28,
    2807 => -28,
    2808 => -28,
    2809 => -29,
    2810 => -29,
    2811 => -29,
    2812 => -29,
    2813 => -29,
    2814 => -29,
    2815 => -29,
    2816 => -29,
    2817 => -29,
    2818 => -29,
    2819 => -29,
    2820 => -29,
    2821 => -29,
    2822 => -29,
    2823 => -29,
    2824 => -29,
    2825 => -29,
    2826 => -29,
    2827 => -29,
    2828 => -29,
    2829 => -29,
    2830 => -29,
    2831 => -29,
    2832 => -29,
    2833 => -29,
    2834 => -29,
    2835 => -29,
    2836 => -29,
    2837 => -29,
    2838 => -29,
    2839 => -29,
    2840 => -29,
    2841 => -29,
    2842 => -29,
    2843 => -29,
    2844 => -29,
    2845 => -29,
    2846 => -29,
    2847 => -29,
    2848 => -29,
    2849 => -29,
    2850 => -29,
    2851 => -29,
    2852 => -29,
    2853 => -29,
    2854 => -29,
    2855 => -29,
    2856 => -29,
    2857 => -29,
    2858 => -29,
    2859 => -29,
    2860 => -29,
    2861 => -29,
    2862 => -29,
    2863 => -29,
    2864 => -29,
    2865 => -29,
    2866 => -29,
    2867 => -29,
    2868 => -29,
    2869 => -30,
    2870 => -30,
    2871 => -30,
    2872 => -30,
    2873 => -30,
    2874 => -30,
    2875 => -30,
    2876 => -30,
    2877 => -30,
    2878 => -30,
    2879 => -30,
    2880 => -30,
    2881 => -30,
    2882 => -30,
    2883 => -30,
    2884 => -30,
    2885 => -30,
    2886 => -30,
    2887 => -30,
    2888 => -30,
    2889 => -30,
    2890 => -30,
    2891 => -30,
    2892 => -30,
    2893 => -30,
    2894 => -30,
    2895 => -30,
    2896 => -30,
    2897 => -30,
    2898 => -30,
    2899 => -30,
    2900 => -30,
    2901 => -30,
    2902 => -30,
    2903 => -30,
    2904 => -30,
    2905 => -30,
    2906 => -30,
    2907 => -30,
    2908 => -30,
    2909 => -30,
    2910 => -30,
    2911 => -30,
    2912 => -30,
    2913 => -30,
    2914 => -30,
    2915 => -30,
    2916 => -30,
    2917 => -30,
    2918 => -30,
    2919 => -30,
    2920 => -30,
    2921 => -30,
    2922 => -30,
    2923 => -30,
    2924 => -30,
    2925 => -30,
    2926 => -30,
    2927 => -30,
    2928 => -30,
    2929 => -30,
    2930 => -30,
    2931 => -30,
    2932 => -30,
    2933 => -30,
    2934 => -30,
    2935 => -30,
    2936 => -30,
    2937 => -30,
    2938 => -30,
    2939 => -30,
    2940 => -30,
    2941 => -30,
    2942 => -30,
    2943 => -30,
    2944 => -30,
    2945 => -30,
    2946 => -30,
    2947 => -30,
    2948 => -30,
    2949 => -30,
    2950 => -30,
    2951 => -30,
    2952 => -30,
    2953 => -30,
    2954 => -30,
    2955 => -31,
    2956 => -31,
    2957 => -31,
    2958 => -31,
    2959 => -31,
    2960 => -31,
    2961 => -31,
    2962 => -31,
    2963 => -31,
    2964 => -31,
    2965 => -31,
    2966 => -31,
    2967 => -31,
    2968 => -31,
    2969 => -31,
    2970 => -31,
    2971 => -31,
    2972 => -31,
    2973 => -31,
    2974 => -31,
    2975 => -31,
    2976 => -31,
    2977 => -31,
    2978 => -31,
    2979 => -31,
    2980 => -31,
    2981 => -31,
    2982 => -31,
    2983 => -31,
    2984 => -31,
    2985 => -31,
    2986 => -31,
    2987 => -31,
    2988 => -31,
    2989 => -31,
    2990 => -31,
    2991 => -31,
    2992 => -31,
    2993 => -31,
    2994 => -31,
    2995 => -31,
    2996 => -31,
    2997 => -31,
    2998 => -31,
    2999 => -31,
    3000 => -31,
    3001 => -31,
    3002 => -31,
    3003 => -31,
    3004 => -31,
    3005 => -31,
    3006 => -31,
    3007 => -31,
    3008 => -31,
    3009 => -31,
    3010 => -31,
    3011 => -31,
    3012 => -31,
    3013 => -31,
    3014 => -31,
    3015 => -31,
    3016 => -31,
    3017 => -31,
    3018 => -31,
    3019 => -31,
    3020 => -31,
    3021 => -31,
    3022 => -31,
    3023 => -31,
    3024 => -31,
    3025 => -31,
    3026 => -31,
    3027 => -31,
    3028 => -31,
    3029 => -31,
    3030 => -31,
    3031 => -31,
    3032 => -31,
    3033 => -31,
    3034 => -31,
    3035 => -31,
    3036 => -31,
    3037 => -31,
    3038 => -31,
    3039 => -31,
    3040 => -31,
    3041 => -31,
    3042 => -31,
    3043 => -31,
    3044 => -31,
    3045 => -31,
    3046 => -31,
    3047 => -31,
    3048 => -31,
    3049 => -31,
    3050 => -31,
    3051 => -31,
    3052 => -31,
    3053 => -31,
    3054 => -31,
    3055 => -31,
    3056 => -31,
    3057 => -31,
    3058 => -31,
    3059 => -31,
    3060 => -31,
    3061 => -31,
    3062 => -31,
    3063 => -31,
    3064 => -31,
    3065 => -31,
    3066 => -31,
    3067 => -31,
    3068 => -31,
    3069 => -31,
    3070 => -31,
    3071 => -31,
    3072 => -31,
    3073 => -31,
    3074 => -31,
    3075 => -31,
    3076 => -31,
    3077 => -31,
    3078 => -31,
    3079 => -31,
    3080 => -31,
    3081 => -31,
    3082 => -31,
    3083 => -31,
    3084 => -31,
    3085 => -31,
    3086 => -31,
    3087 => -31,
    3088 => -31,
    3089 => -31,
    3090 => -31,
    3091 => -31,
    3092 => -31,
    3093 => -31,
    3094 => -31,
    3095 => -31,
    3096 => -31,
    3097 => -31,
    3098 => -31,
    3099 => -31,
    3100 => -31,
    3101 => -31,
    3102 => -31,
    3103 => -31,
    3104 => -31,
    3105 => -31,
    3106 => -31,
    3107 => -31,
    3108 => -31,
    3109 => -31,
    3110 => -31,
    3111 => -31,
    3112 => -31,
    3113 => -31,
    3114 => -31,
    3115 => -31,
    3116 => -31,
    3117 => -31,
    3118 => -31,
    3119 => -31,
    3120 => -31,
    3121 => -31,
    3122 => -31,
    3123 => -31,
    3124 => -31,
    3125 => -31,
    3126 => -31,
    3127 => -31,
    3128 => -31,
    3129 => -31,
    3130 => -31,
    3131 => -31,
    3132 => -31,
    3133 => -31,
    3134 => -31,
    3135 => -31,
    3136 => -31,
    3137 => -31,
    3138 => -31,
    3139 => -31,
    3140 => -31,
    3141 => -31,
    3142 => -31,
    3143 => -31,
    3144 => -31,
    3145 => -31,
    3146 => -31,
    3147 => -31,
    3148 => -31,
    3149 => -31,
    3150 => -31,
    3151 => -31,
    3152 => -31,
    3153 => -31,
    3154 => -31,
    3155 => -31,
    3156 => -31,
    3157 => -31,
    3158 => -31,
    3159 => -31,
    3160 => -31,
    3161 => -31,
    3162 => -31,
    3163 => -31,
    3164 => -31,
    3165 => -31,
    3166 => -31,
    3167 => -31,
    3168 => -31,
    3169 => -31,
    3170 => -31,
    3171 => -31,
    3172 => -31,
    3173 => -31,
    3174 => -31,
    3175 => -31,
    3176 => -31,
    3177 => -31,
    3178 => -31,
    3179 => -31,
    3180 => -31,
    3181 => -31,
    3182 => -31,
    3183 => -31,
    3184 => -31,
    3185 => -31,
    3186 => -31,
    3187 => -31,
    3188 => -31,
    3189 => -31,
    3190 => -30,
    3191 => -30,
    3192 => -30,
    3193 => -30,
    3194 => -30,
    3195 => -30,
    3196 => -30,
    3197 => -30,
    3198 => -30,
    3199 => -30,
    3200 => -30,
    3201 => -30,
    3202 => -30,
    3203 => -30,
    3204 => -30,
    3205 => -30,
    3206 => -30,
    3207 => -30,
    3208 => -30,
    3209 => -30,
    3210 => -30,
    3211 => -30,
    3212 => -30,
    3213 => -30,
    3214 => -30,
    3215 => -30,
    3216 => -30,
    3217 => -30,
    3218 => -30,
    3219 => -30,
    3220 => -30,
    3221 => -30,
    3222 => -30,
    3223 => -30,
    3224 => -30,
    3225 => -30,
    3226 => -30,
    3227 => -30,
    3228 => -30,
    3229 => -30,
    3230 => -30,
    3231 => -30,
    3232 => -30,
    3233 => -30,
    3234 => -30,
    3235 => -30,
    3236 => -30,
    3237 => -30,
    3238 => -30,
    3239 => -30,
    3240 => -30,
    3241 => -30,
    3242 => -30,
    3243 => -30,
    3244 => -30,
    3245 => -30,
    3246 => -30,
    3247 => -30,
    3248 => -30,
    3249 => -30,
    3250 => -30,
    3251 => -30,
    3252 => -30,
    3253 => -30,
    3254 => -30,
    3255 => -30,
    3256 => -30,
    3257 => -30,
    3258 => -30,
    3259 => -30,
    3260 => -30,
    3261 => -30,
    3262 => -30,
    3263 => -30,
    3264 => -30,
    3265 => -30,
    3266 => -30,
    3267 => -30,
    3268 => -30,
    3269 => -30,
    3270 => -30,
    3271 => -30,
    3272 => -30,
    3273 => -30,
    3274 => -30,
    3275 => -30,
    3276 => -29,
    3277 => -29,
    3278 => -29,
    3279 => -29,
    3280 => -29,
    3281 => -29,
    3282 => -29,
    3283 => -29,
    3284 => -29,
    3285 => -29,
    3286 => -29,
    3287 => -29,
    3288 => -29,
    3289 => -29,
    3290 => -29,
    3291 => -29,
    3292 => -29,
    3293 => -29,
    3294 => -29,
    3295 => -29,
    3296 => -29,
    3297 => -29,
    3298 => -29,
    3299 => -29,
    3300 => -29,
    3301 => -29,
    3302 => -29,
    3303 => -29,
    3304 => -29,
    3305 => -29,
    3306 => -29,
    3307 => -29,
    3308 => -29,
    3309 => -29,
    3310 => -29,
    3311 => -29,
    3312 => -29,
    3313 => -29,
    3314 => -29,
    3315 => -29,
    3316 => -29,
    3317 => -29,
    3318 => -29,
    3319 => -29,
    3320 => -29,
    3321 => -29,
    3322 => -29,
    3323 => -29,
    3324 => -29,
    3325 => -29,
    3326 => -29,
    3327 => -29,
    3328 => -29,
    3329 => -29,
    3330 => -29,
    3331 => -29,
    3332 => -29,
    3333 => -29,
    3334 => -29,
    3335 => -29,
    3336 => -28,
    3337 => -28,
    3338 => -28,
    3339 => -28,
    3340 => -28,
    3341 => -28,
    3342 => -28,
    3343 => -28,
    3344 => -28,
    3345 => -28,
    3346 => -28,
    3347 => -28,
    3348 => -28,
    3349 => -28,
    3350 => -28,
    3351 => -28,
    3352 => -28,
    3353 => -28,
    3354 => -28,
    3355 => -28,
    3356 => -28,
    3357 => -28,
    3358 => -28,
    3359 => -28,
    3360 => -28,
    3361 => -28,
    3362 => -28,
    3363 => -28,
    3364 => -28,
    3365 => -28,
    3366 => -28,
    3367 => -28,
    3368 => -28,
    3369 => -28,
    3370 => -28,
    3371 => -28,
    3372 => -28,
    3373 => -28,
    3374 => -28,
    3375 => -28,
    3376 => -28,
    3377 => -28,
    3378 => -28,
    3379 => -28,
    3380 => -28,
    3381 => -28,
    3382 => -28,
    3383 => -28,
    3384 => -28,
    3385 => -27,
    3386 => -27,
    3387 => -27,
    3388 => -27,
    3389 => -27,
    3390 => -27,
    3391 => -27,
    3392 => -27,
    3393 => -27,
    3394 => -27,
    3395 => -27,
    3396 => -27,
    3397 => -27,
    3398 => -27,
    3399 => -27,
    3400 => -27,
    3401 => -27,
    3402 => -27,
    3403 => -27,
    3404 => -27,
    3405 => -27,
    3406 => -27,
    3407 => -27,
    3408 => -27,
    3409 => -27,
    3410 => -27,
    3411 => -27,
    3412 => -27,
    3413 => -27,
    3414 => -27,
    3415 => -27,
    3416 => -27,
    3417 => -27,
    3418 => -27,
    3419 => -27,
    3420 => -27,
    3421 => -27,
    3422 => -27,
    3423 => -27,
    3424 => -27,
    3425 => -27,
    3426 => -27,
    3427 => -27,
    3428 => -26,
    3429 => -26,
    3430 => -26,
    3431 => -26,
    3432 => -26,
    3433 => -26,
    3434 => -26,
    3435 => -26,
    3436 => -26,
    3437 => -26,
    3438 => -26,
    3439 => -26,
    3440 => -26,
    3441 => -26,
    3442 => -26,
    3443 => -26,
    3444 => -26,
    3445 => -26,
    3446 => -26,
    3447 => -26,
    3448 => -26,
    3449 => -26,
    3450 => -26,
    3451 => -26,
    3452 => -26,
    3453 => -26,
    3454 => -26,
    3455 => -26,
    3456 => -26,
    3457 => -26,
    3458 => -26,
    3459 => -26,
    3460 => -26,
    3461 => -26,
    3462 => -26,
    3463 => -26,
    3464 => -26,
    3465 => -26,
    3466 => -26,
    3467 => -25,
    3468 => -25,
    3469 => -25,
    3470 => -25,
    3471 => -25,
    3472 => -25,
    3473 => -25,
    3474 => -25,
    3475 => -25,
    3476 => -25,
    3477 => -25,
    3478 => -25,
    3479 => -25,
    3480 => -25,
    3481 => -25,
    3482 => -25,
    3483 => -25,
    3484 => -25,
    3485 => -25,
    3486 => -25,
    3487 => -25,
    3488 => -25,
    3489 => -25,
    3490 => -25,
    3491 => -25,
    3492 => -25,
    3493 => -25,
    3494 => -25,
    3495 => -25,
    3496 => -25,
    3497 => -25,
    3498 => -25,
    3499 => -25,
    3500 => -25,
    3501 => -25,
    3502 => -24,
    3503 => -24,
    3504 => -24,
    3505 => -24,
    3506 => -24,
    3507 => -24,
    3508 => -24,
    3509 => -24,
    3510 => -24,
    3511 => -24,
    3512 => -24,
    3513 => -24,
    3514 => -24,
    3515 => -24,
    3516 => -24,
    3517 => -24,
    3518 => -24,
    3519 => -24,
    3520 => -24,
    3521 => -24,
    3522 => -24,
    3523 => -24,
    3524 => -24,
    3525 => -24,
    3526 => -24,
    3527 => -24,
    3528 => -24,
    3529 => -24,
    3530 => -24,
    3531 => -24,
    3532 => -24,
    3533 => -24,
    3534 => -24,
    3535 => -24,
    3536 => -23,
    3537 => -23,
    3538 => -23,
    3539 => -23,
    3540 => -23,
    3541 => -23,
    3542 => -23,
    3543 => -23,
    3544 => -23,
    3545 => -23,
    3546 => -23,
    3547 => -23,
    3548 => -23,
    3549 => -23,
    3550 => -23,
    3551 => -23,
    3552 => -23,
    3553 => -23,
    3554 => -23,
    3555 => -23,
    3556 => -23,
    3557 => -23,
    3558 => -23,
    3559 => -23,
    3560 => -23,
    3561 => -23,
    3562 => -23,
    3563 => -23,
    3564 => -23,
    3565 => -23,
    3566 => -23,
    3567 => -22,
    3568 => -22,
    3569 => -22,
    3570 => -22,
    3571 => -22,
    3572 => -22,
    3573 => -22,
    3574 => -22,
    3575 => -22,
    3576 => -22,
    3577 => -22,
    3578 => -22,
    3579 => -22,
    3580 => -22,
    3581 => -22,
    3582 => -22,
    3583 => -22,
    3584 => -22,
    3585 => -22,
    3586 => -22,
    3587 => -22,
    3588 => -22,
    3589 => -22,
    3590 => -22,
    3591 => -22,
    3592 => -22,
    3593 => -22,
    3594 => -22,
    3595 => -22,
    3596 => -22,
    3597 => -21,
    3598 => -21,
    3599 => -21,
    3600 => -21,
    3601 => -21,
    3602 => -21,
    3603 => -21,
    3604 => -21,
    3605 => -21,
    3606 => -21,
    3607 => -21,
    3608 => -21,
    3609 => -21,
    3610 => -21,
    3611 => -21,
    3612 => -21,
    3613 => -21,
    3614 => -21,
    3615 => -21,
    3616 => -21,
    3617 => -21,
    3618 => -21,
    3619 => -21,
    3620 => -21,
    3621 => -21,
    3622 => -21,
    3623 => -21,
    3624 => -21,
    3625 => -20,
    3626 => -20,
    3627 => -20,
    3628 => -20,
    3629 => -20,
    3630 => -20,
    3631 => -20,
    3632 => -20,
    3633 => -20,
    3634 => -20,
    3635 => -20,
    3636 => -20,
    3637 => -20,
    3638 => -20,
    3639 => -20,
    3640 => -20,
    3641 => -20,
    3642 => -20,
    3643 => -20,
    3644 => -20,
    3645 => -20,
    3646 => -20,
    3647 => -20,
    3648 => -20,
    3649 => -20,
    3650 => -20,
    3651 => -20,
    3652 => -20,
    3653 => -19,
    3654 => -19,
    3655 => -19,
    3656 => -19,
    3657 => -19,
    3658 => -19,
    3659 => -19,
    3660 => -19,
    3661 => -19,
    3662 => -19,
    3663 => -19,
    3664 => -19,
    3665 => -19,
    3666 => -19,
    3667 => -19,
    3668 => -19,
    3669 => -19,
    3670 => -19,
    3671 => -19,
    3672 => -19,
    3673 => -19,
    3674 => -19,
    3675 => -19,
    3676 => -19,
    3677 => -19,
    3678 => -19,
    3679 => -19,
    3680 => -18,
    3681 => -18,
    3682 => -18,
    3683 => -18,
    3684 => -18,
    3685 => -18,
    3686 => -18,
    3687 => -18,
    3688 => -18,
    3689 => -18,
    3690 => -18,
    3691 => -18,
    3692 => -18,
    3693 => -18,
    3694 => -18,
    3695 => -18,
    3696 => -18,
    3697 => -18,
    3698 => -18,
    3699 => -18,
    3700 => -18,
    3701 => -18,
    3702 => -18,
    3703 => -18,
    3704 => -18,
    3705 => -17,
    3706 => -17,
    3707 => -17,
    3708 => -17,
    3709 => -17,
    3710 => -17,
    3711 => -17,
    3712 => -17,
    3713 => -17,
    3714 => -17,
    3715 => -17,
    3716 => -17,
    3717 => -17,
    3718 => -17,
    3719 => -17,
    3720 => -17,
    3721 => -17,
    3722 => -17,
    3723 => -17,
    3724 => -17,
    3725 => -17,
    3726 => -17,
    3727 => -17,
    3728 => -17,
    3729 => -17,
    3730 => -17,
    3731 => -16,
    3732 => -16,
    3733 => -16,
    3734 => -16,
    3735 => -16,
    3736 => -16,
    3737 => -16,
    3738 => -16,
    3739 => -16,
    3740 => -16,
    3741 => -16,
    3742 => -16,
    3743 => -16,
    3744 => -16,
    3745 => -16,
    3746 => -16,
    3747 => -16,
    3748 => -16,
    3749 => -16,
    3750 => -16,
    3751 => -16,
    3752 => -16,
    3753 => -16,
    3754 => -16,
    3755 => -15,
    3756 => -15,
    3757 => -15,
    3758 => -15,
    3759 => -15,
    3760 => -15,
    3761 => -15,
    3762 => -15,
    3763 => -15,
    3764 => -15,
    3765 => -15,
    3766 => -15,
    3767 => -15,
    3768 => -15,
    3769 => -15,
    3770 => -15,
    3771 => -15,
    3772 => -15,
    3773 => -15,
    3774 => -15,
    3775 => -15,
    3776 => -15,
    3777 => -15,
    3778 => -15,
    3779 => -14,
    3780 => -14,
    3781 => -14,
    3782 => -14,
    3783 => -14,
    3784 => -14,
    3785 => -14,
    3786 => -14,
    3787 => -14,
    3788 => -14,
    3789 => -14,
    3790 => -14,
    3791 => -14,
    3792 => -14,
    3793 => -14,
    3794 => -14,
    3795 => -14,
    3796 => -14,
    3797 => -14,
    3798 => -14,
    3799 => -14,
    3800 => -14,
    3801 => -14,
    3802 => -14,
    3803 => -13,
    3804 => -13,
    3805 => -13,
    3806 => -13,
    3807 => -13,
    3808 => -13,
    3809 => -13,
    3810 => -13,
    3811 => -13,
    3812 => -13,
    3813 => -13,
    3814 => -13,
    3815 => -13,
    3816 => -13,
    3817 => -13,
    3818 => -13,
    3819 => -13,
    3820 => -13,
    3821 => -13,
    3822 => -13,
    3823 => -13,
    3824 => -13,
    3825 => -13,
    3826 => -12,
    3827 => -12,
    3828 => -12,
    3829 => -12,
    3830 => -12,
    3831 => -12,
    3832 => -12,
    3833 => -12,
    3834 => -12,
    3835 => -12,
    3836 => -12,
    3837 => -12,
    3838 => -12,
    3839 => -12,
    3840 => -12,
    3841 => -12,
    3842 => -12,
    3843 => -12,
    3844 => -12,
    3845 => -12,
    3846 => -12,
    3847 => -12,
    3848 => -12,
    3849 => -11,
    3850 => -11,
    3851 => -11,
    3852 => -11,
    3853 => -11,
    3854 => -11,
    3855 => -11,
    3856 => -11,
    3857 => -11,
    3858 => -11,
    3859 => -11,
    3860 => -11,
    3861 => -11,
    3862 => -11,
    3863 => -11,
    3864 => -11,
    3865 => -11,
    3866 => -11,
    3867 => -11,
    3868 => -11,
    3869 => -11,
    3870 => -11,
    3871 => -10,
    3872 => -10,
    3873 => -10,
    3874 => -10,
    3875 => -10,
    3876 => -10,
    3877 => -10,
    3878 => -10,
    3879 => -10,
    3880 => -10,
    3881 => -10,
    3882 => -10,
    3883 => -10,
    3884 => -10,
    3885 => -10,
    3886 => -10,
    3887 => -10,
    3888 => -10,
    3889 => -10,
    3890 => -10,
    3891 => -10,
    3892 => -10,
    3893 => -9,
    3894 => -9,
    3895 => -9,
    3896 => -9,
    3897 => -9,
    3898 => -9,
    3899 => -9,
    3900 => -9,
    3901 => -9,
    3902 => -9,
    3903 => -9,
    3904 => -9,
    3905 => -9,
    3906 => -9,
    3907 => -9,
    3908 => -9,
    3909 => -9,
    3910 => -9,
    3911 => -9,
    3912 => -9,
    3913 => -9,
    3914 => -9,
    3915 => -8,
    3916 => -8,
    3917 => -8,
    3918 => -8,
    3919 => -8,
    3920 => -8,
    3921 => -8,
    3922 => -8,
    3923 => -8,
    3924 => -8,
    3925 => -8,
    3926 => -8,
    3927 => -8,
    3928 => -8,
    3929 => -8,
    3930 => -8,
    3931 => -8,
    3932 => -8,
    3933 => -8,
    3934 => -8,
    3935 => -8,
    3936 => -8,
    3937 => -7,
    3938 => -7,
    3939 => -7,
    3940 => -7,
    3941 => -7,
    3942 => -7,
    3943 => -7,
    3944 => -7,
    3945 => -7,
    3946 => -7,
    3947 => -7,
    3948 => -7,
    3949 => -7,
    3950 => -7,
    3951 => -7,
    3952 => -7,
    3953 => -7,
    3954 => -7,
    3955 => -7,
    3956 => -7,
    3957 => -7,
    3958 => -7,
    3959 => -6,
    3960 => -6,
    3961 => -6,
    3962 => -6,
    3963 => -6,
    3964 => -6,
    3965 => -6,
    3966 => -6,
    3967 => -6,
    3968 => -6,
    3969 => -6,
    3970 => -6,
    3971 => -6,
    3972 => -6,
    3973 => -6,
    3974 => -6,
    3975 => -6,
    3976 => -6,
    3977 => -6,
    3978 => -6,
    3979 => -6,
    3980 => -5,
    3981 => -5,
    3982 => -5,
    3983 => -5,
    3984 => -5,
    3985 => -5,
    3986 => -5,
    3987 => -5,
    3988 => -5,
    3989 => -5,
    3990 => -5,
    3991 => -5,
    3992 => -5,
    3993 => -5,
    3994 => -5,
    3995 => -5,
    3996 => -5,
    3997 => -5,
    3998 => -5,
    3999 => -5,
    4000 => -5,
    4001 => -5,
    4002 => -4,
    4003 => -4,
    4004 => -4,
    4005 => -4,
    4006 => -4,
    4007 => -4,
    4008 => -4,
    4009 => -4,
    4010 => -4,
    4011 => -4,
    4012 => -4,
    4013 => -4,
    4014 => -4,
    4015 => -4,
    4016 => -4,
    4017 => -4,
    4018 => -4,
    4019 => -4,
    4020 => -4,
    4021 => -4,
    4022 => -4,
    4023 => -3,
    4024 => -3,
    4025 => -3,
    4026 => -3,
    4027 => -3,
    4028 => -3,
    4029 => -3,
    4030 => -3,
    4031 => -3,
    4032 => -3,
    4033 => -3,
    4034 => -3,
    4035 => -3,
    4036 => -3,
    4037 => -3,
    4038 => -3,
    4039 => -3,
    4040 => -3,
    4041 => -3,
    4042 => -3,
    4043 => -3,
    4044 => -2,
    4045 => -2,
    4046 => -2,
    4047 => -2,
    4048 => -2,
    4049 => -2,
    4050 => -2,
    4051 => -2,
    4052 => -2,
    4053 => -2,
    4054 => -2,
    4055 => -2,
    4056 => -2,
    4057 => -2,
    4058 => -2,
    4059 => -2,
    4060 => -2,
    4061 => -2,
    4062 => -2,
    4063 => -2,
    4064 => -2,
    4065 => -1,
    4066 => -1,
    4067 => -1,
    4068 => -1,
    4069 => -1,
    4070 => -1,
    4071 => -1,
    4072 => -1,
    4073 => -1,
    4074 => -1,
    4075 => -1,
    4076 => -1,
    4077 => -1,
    4078 => -1,
    4079 => -1,
    4080 => -1,
    4081 => -1,
    4082 => -1,
    4083 => -1,
    4084 => -1,
    4085 => -1,
    4086 => 0,
    4087 => 0,
    4088 => 0,
    4089 => 0,
    4090 => 0,
    4091 => 0,
    4092 => 0,
    4093 => 0,
    4094 => 0,
    4095 => 0
  );

begin
  ddfs_out <= std_logic_vector(to_signed(LUT(to_integer(unsigned(address))),6));
end architecture;

library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity ddfs_qlut_1024_6bit is
  port (
    address  : in  std_logic_vector(9 downto 0);
    ddfs_out : out std_logic_vector(5 downto 0)
  );
end entity;

architecture rtl of ddfs_qlut_1024_6bit is

  type LUT_t is array (natural range 0 to 1023) of integer;
  constant LUT: LUT_t := (
    0 => 0,
    1 => 0,
    2 => 0,
    3 => 0,
    4 => 0,
    5 => 0,
    6 => 0,
    7 => 0,
    8 => 0,
    9 => 0,
    10 => 0,
    11 => 1,
    12 => 1,
    13 => 1,
    14 => 1,
    15 => 1,
    16 => 1,
    17 => 1,
    18 => 1,
    19 => 1,
    20 => 1,
    21 => 1,
    22 => 1,
    23 => 1,
    24 => 1,
    25 => 1,
    26 => 1,
    27 => 1,
    28 => 1,
    29 => 1,
    30 => 1,
    31 => 1,
    32 => 2,
    33 => 2,
    34 => 2,
    35 => 2,
    36 => 2,
    37 => 2,
    38 => 2,
    39 => 2,
    40 => 2,
    41 => 2,
    42 => 2,
    43 => 2,
    44 => 2,
    45 => 2,
    46 => 2,
    47 => 2,
    48 => 2,
    49 => 2,
    50 => 2,
    51 => 2,
    52 => 2,
    53 => 3,
    54 => 3,
    55 => 3,
    56 => 3,
    57 => 3,
    58 => 3,
    59 => 3,
    60 => 3,
    61 => 3,
    62 => 3,
    63 => 3,
    64 => 3,
    65 => 3,
    66 => 3,
    67 => 3,
    68 => 3,
    69 => 3,
    70 => 3,
    71 => 3,
    72 => 3,
    73 => 3,
    74 => 4,
    75 => 4,
    76 => 4,
    77 => 4,
    78 => 4,
    79 => 4,
    80 => 4,
    81 => 4,
    82 => 4,
    83 => 4,
    84 => 4,
    85 => 4,
    86 => 4,
    87 => 4,
    88 => 4,
    89 => 4,
    90 => 4,
    91 => 4,
    92 => 4,
    93 => 4,
    94 => 4,
    95 => 5,
    96 => 5,
    97 => 5,
    98 => 5,
    99 => 5,
    100 => 5,
    101 => 5,
    102 => 5,
    103 => 5,
    104 => 5,
    105 => 5,
    106 => 5,
    107 => 5,
    108 => 5,
    109 => 5,
    110 => 5,
    111 => 5,
    112 => 5,
    113 => 5,
    114 => 5,
    115 => 5,
    116 => 5,
    117 => 6,
    118 => 6,
    119 => 6,
    120 => 6,
    121 => 6,
    122 => 6,
    123 => 6,
    124 => 6,
    125 => 6,
    126 => 6,
    127 => 6,
    128 => 6,
    129 => 6,
    130 => 6,
    131 => 6,
    132 => 6,
    133 => 6,
    134 => 6,
    135 => 6,
    136 => 6,
    137 => 6,
    138 => 7,
    139 => 7,
    140 => 7,
    141 => 7,
    142 => 7,
    143 => 7,
    144 => 7,
    145 => 7,
    146 => 7,
    147 => 7,
    148 => 7,
    149 => 7,
    150 => 7,
    151 => 7,
    152 => 7,
    153 => 7,
    154 => 7,
    155 => 7,
    156 => 7,
    157 => 7,
    158 => 7,
    159 => 7,
    160 => 8,
    161 => 8,
    162 => 8,
    163 => 8,
    164 => 8,
    165 => 8,
    166 => 8,
    167 => 8,
    168 => 8,
    169 => 8,
    170 => 8,
    171 => 8,
    172 => 8,
    173 => 8,
    174 => 8,
    175 => 8,
    176 => 8,
    177 => 8,
    178 => 8,
    179 => 8,
    180 => 8,
    181 => 8,
    182 => 9,
    183 => 9,
    184 => 9,
    185 => 9,
    186 => 9,
    187 => 9,
    188 => 9,
    189 => 9,
    190 => 9,
    191 => 9,
    192 => 9,
    193 => 9,
    194 => 9,
    195 => 9,
    196 => 9,
    197 => 9,
    198 => 9,
    199 => 9,
    200 => 9,
    201 => 9,
    202 => 9,
    203 => 9,
    204 => 10,
    205 => 10,
    206 => 10,
    207 => 10,
    208 => 10,
    209 => 10,
    210 => 10,
    211 => 10,
    212 => 10,
    213 => 10,
    214 => 10,
    215 => 10,
    216 => 10,
    217 => 10,
    218 => 10,
    219 => 10,
    220 => 10,
    221 => 10,
    222 => 10,
    223 => 10,
    224 => 10,
    225 => 10,
    226 => 11,
    227 => 11,
    228 => 11,
    229 => 11,
    230 => 11,
    231 => 11,
    232 => 11,
    233 => 11,
    234 => 11,
    235 => 11,
    236 => 11,
    237 => 11,
    238 => 11,
    239 => 11,
    240 => 11,
    241 => 11,
    242 => 11,
    243 => 11,
    244 => 11,
    245 => 11,
    246 => 11,
    247 => 11,
    248 => 12,
    249 => 12,
    250 => 12,
    251 => 12,
    252 => 12,
    253 => 12,
    254 => 12,
    255 => 12,
    256 => 12,
    257 => 12,
    258 => 12,
    259 => 12,
    260 => 12,
    261 => 12,
    262 => 12,
    263 => 12,
    264 => 12,
    265 => 12,
    266 => 12,
    267 => 12,
    268 => 12,
    269 => 12,
    270 => 12,
    271 => 13,
    272 => 13,
    273 => 13,
    274 => 13,
    275 => 13,
    276 => 13,
    277 => 13,
    278 => 13,
    279 => 13,
    280 => 13,
    281 => 13,
    282 => 13,
    283 => 13,
    284 => 13,
    285 => 13,
    286 => 13,
    287 => 13,
    288 => 13,
    289 => 13,
    290 => 13,
    291 => 13,
    292 => 13,
    293 => 13,
    294 => 14,
    295 => 14,
    296 => 14,
    297 => 14,
    298 => 14,
    299 => 14,
    300 => 14,
    301 => 14,
    302 => 14,
    303 => 14,
    304 => 14,
    305 => 14,
    306 => 14,
    307 => 14,
    308 => 14,
    309 => 14,
    310 => 14,
    311 => 14,
    312 => 14,
    313 => 14,
    314 => 14,
    315 => 14,
    316 => 14,
    317 => 14,
    318 => 15,
    319 => 15,
    320 => 15,
    321 => 15,
    322 => 15,
    323 => 15,
    324 => 15,
    325 => 15,
    326 => 15,
    327 => 15,
    328 => 15,
    329 => 15,
    330 => 15,
    331 => 15,
    332 => 15,
    333 => 15,
    334 => 15,
    335 => 15,
    336 => 15,
    337 => 15,
    338 => 15,
    339 => 15,
    340 => 15,
    341 => 15,
    342 => 16,
    343 => 16,
    344 => 16,
    345 => 16,
    346 => 16,
    347 => 16,
    348 => 16,
    349 => 16,
    350 => 16,
    351 => 16,
    352 => 16,
    353 => 16,
    354 => 16,
    355 => 16,
    356 => 16,
    357 => 16,
    358 => 16,
    359 => 16,
    360 => 16,
    361 => 16,
    362 => 16,
    363 => 16,
    364 => 16,
    365 => 16,
    366 => 17,
    367 => 17,
    368 => 17,
    369 => 17,
    370 => 17,
    371 => 17,
    372 => 17,
    373 => 17,
    374 => 17,
    375 => 17,
    376 => 17,
    377 => 17,
    378 => 17,
    379 => 17,
    380 => 17,
    381 => 17,
    382 => 17,
    383 => 17,
    384 => 17,
    385 => 17,
    386 => 17,
    387 => 17,
    388 => 17,
    389 => 17,
    390 => 17,
    391 => 17,
    392 => 18,
    393 => 18,
    394 => 18,
    395 => 18,
    396 => 18,
    397 => 18,
    398 => 18,
    399 => 18,
    400 => 18,
    401 => 18,
    402 => 18,
    403 => 18,
    404 => 18,
    405 => 18,
    406 => 18,
    407 => 18,
    408 => 18,
    409 => 18,
    410 => 18,
    411 => 18,
    412 => 18,
    413 => 18,
    414 => 18,
    415 => 18,
    416 => 18,
    417 => 19,
    418 => 19,
    419 => 19,
    420 => 19,
    421 => 19,
    422 => 19,
    423 => 19,
    424 => 19,
    425 => 19,
    426 => 19,
    427 => 19,
    428 => 19,
    429 => 19,
    430 => 19,
    431 => 19,
    432 => 19,
    433 => 19,
    434 => 19,
    435 => 19,
    436 => 19,
    437 => 19,
    438 => 19,
    439 => 19,
    440 => 19,
    441 => 19,
    442 => 19,
    443 => 19,
    444 => 20,
    445 => 20,
    446 => 20,
    447 => 20,
    448 => 20,
    449 => 20,
    450 => 20,
    451 => 20,
    452 => 20,
    453 => 20,
    454 => 20,
    455 => 20,
    456 => 20,
    457 => 20,
    458 => 20,
    459 => 20,
    460 => 20,
    461 => 20,
    462 => 20,
    463 => 20,
    464 => 20,
    465 => 20,
    466 => 20,
    467 => 20,
    468 => 20,
    469 => 20,
    470 => 20,
    471 => 20,
    472 => 21,
    473 => 21,
    474 => 21,
    475 => 21,
    476 => 21,
    477 => 21,
    478 => 21,
    479 => 21,
    480 => 21,
    481 => 21,
    482 => 21,
    483 => 21,
    484 => 21,
    485 => 21,
    486 => 21,
    487 => 21,
    488 => 21,
    489 => 21,
    490 => 21,
    491 => 21,
    492 => 21,
    493 => 21,
    494 => 21,
    495 => 21,
    496 => 21,
    497 => 21,
    498 => 21,
    499 => 21,
    500 => 22,
    501 => 22,
    502 => 22,
    503 => 22,
    504 => 22,
    505 => 22,
    506 => 22,
    507 => 22,
    508 => 22,
    509 => 22,
    510 => 22,
    511 => 22,
    512 => 22,
    513 => 22,
    514 => 22,
    515 => 22,
    516 => 22,
    517 => 22,
    518 => 22,
    519 => 22,
    520 => 22,
    521 => 22,
    522 => 22,
    523 => 22,
    524 => 22,
    525 => 22,
    526 => 22,
    527 => 22,
    528 => 22,
    529 => 22,
    530 => 23,
    531 => 23,
    532 => 23,
    533 => 23,
    534 => 23,
    535 => 23,
    536 => 23,
    537 => 23,
    538 => 23,
    539 => 23,
    540 => 23,
    541 => 23,
    542 => 23,
    543 => 23,
    544 => 23,
    545 => 23,
    546 => 23,
    547 => 23,
    548 => 23,
    549 => 23,
    550 => 23,
    551 => 23,
    552 => 23,
    553 => 23,
    554 => 23,
    555 => 23,
    556 => 23,
    557 => 23,
    558 => 23,
    559 => 23,
    560 => 23,
    561 => 24,
    562 => 24,
    563 => 24,
    564 => 24,
    565 => 24,
    566 => 24,
    567 => 24,
    568 => 24,
    569 => 24,
    570 => 24,
    571 => 24,
    572 => 24,
    573 => 24,
    574 => 24,
    575 => 24,
    576 => 24,
    577 => 24,
    578 => 24,
    579 => 24,
    580 => 24,
    581 => 24,
    582 => 24,
    583 => 24,
    584 => 24,
    585 => 24,
    586 => 24,
    587 => 24,
    588 => 24,
    589 => 24,
    590 => 24,
    591 => 24,
    592 => 24,
    593 => 24,
    594 => 24,
    595 => 25,
    596 => 25,
    597 => 25,
    598 => 25,
    599 => 25,
    600 => 25,
    601 => 25,
    602 => 25,
    603 => 25,
    604 => 25,
    605 => 25,
    606 => 25,
    607 => 25,
    608 => 25,
    609 => 25,
    610 => 25,
    611 => 25,
    612 => 25,
    613 => 25,
    614 => 25,
    615 => 25,
    616 => 25,
    617 => 25,
    618 => 25,
    619 => 25,
    620 => 25,
    621 => 25,
    622 => 25,
    623 => 25,
    624 => 25,
    625 => 25,
    626 => 25,
    627 => 25,
    628 => 25,
    629 => 25,
    630 => 26,
    631 => 26,
    632 => 26,
    633 => 26,
    634 => 26,
    635 => 26,
    636 => 26,
    637 => 26,
    638 => 26,
    639 => 26,
    640 => 26,
    641 => 26,
    642 => 26,
    643 => 26,
    644 => 26,
    645 => 26,
    646 => 26,
    647 => 26,
    648 => 26,
    649 => 26,
    650 => 26,
    651 => 26,
    652 => 26,
    653 => 26,
    654 => 26,
    655 => 26,
    656 => 26,
    657 => 26,
    658 => 26,
    659 => 26,
    660 => 26,
    661 => 26,
    662 => 26,
    663 => 26,
    664 => 26,
    665 => 26,
    666 => 26,
    667 => 26,
    668 => 26,
    669 => 27,
    670 => 27,
    671 => 27,
    672 => 27,
    673 => 27,
    674 => 27,
    675 => 27,
    676 => 27,
    677 => 27,
    678 => 27,
    679 => 27,
    680 => 27,
    681 => 27,
    682 => 27,
    683 => 27,
    684 => 27,
    685 => 27,
    686 => 27,
    687 => 27,
    688 => 27,
    689 => 27,
    690 => 27,
    691 => 27,
    692 => 27,
    693 => 27,
    694 => 27,
    695 => 27,
    696 => 27,
    697 => 27,
    698 => 27,
    699 => 27,
    700 => 27,
    701 => 27,
    702 => 27,
    703 => 27,
    704 => 27,
    705 => 27,
    706 => 27,
    707 => 27,
    708 => 27,
    709 => 27,
    710 => 27,
    711 => 27,
    712 => 28,
    713 => 28,
    714 => 28,
    715 => 28,
    716 => 28,
    717 => 28,
    718 => 28,
    719 => 28,
    720 => 28,
    721 => 28,
    722 => 28,
    723 => 28,
    724 => 28,
    725 => 28,
    726 => 28,
    727 => 28,
    728 => 28,
    729 => 28,
    730 => 28,
    731 => 28,
    732 => 28,
    733 => 28,
    734 => 28,
    735 => 28,
    736 => 28,
    737 => 28,
    738 => 28,
    739 => 28,
    740 => 28,
    741 => 28,
    742 => 28,
    743 => 28,
    744 => 28,
    745 => 28,
    746 => 28,
    747 => 28,
    748 => 28,
    749 => 28,
    750 => 28,
    751 => 28,
    752 => 28,
    753 => 28,
    754 => 28,
    755 => 28,
    756 => 28,
    757 => 28,
    758 => 28,
    759 => 28,
    760 => 28,
    761 => 29,
    762 => 29,
    763 => 29,
    764 => 29,
    765 => 29,
    766 => 29,
    767 => 29,
    768 => 29,
    769 => 29,
    770 => 29,
    771 => 29,
    772 => 29,
    773 => 29,
    774 => 29,
    775 => 29,
    776 => 29,
    777 => 29,
    778 => 29,
    779 => 29,
    780 => 29,
    781 => 29,
    782 => 29,
    783 => 29,
    784 => 29,
    785 => 29,
    786 => 29,
    787 => 29,
    788 => 29,
    789 => 29,
    790 => 29,
    791 => 29,
    792 => 29,
    793 => 29,
    794 => 29,
    795 => 29,
    796 => 29,
    797 => 29,
    798 => 29,
    799 => 29,
    800 => 29,
    801 => 29,
    802 => 29,
    803 => 29,
    804 => 29,
    805 => 29,
    806 => 29,
    807 => 29,
    808 => 29,
    809 => 29,
    810 => 29,
    811 => 29,
    812 => 29,
    813 => 29,
    814 => 29,
    815 => 29,
    816 => 29,
    817 => 29,
    818 => 29,
    819 => 29,
    820 => 29,
    821 => 30,
    822 => 30,
    823 => 30,
    824 => 30,
    825 => 30,
    826 => 30,
    827 => 30,
    828 => 30,
    829 => 30,
    830 => 30,
    831 => 30,
    832 => 30,
    833 => 30,
    834 => 30,
    835 => 30,
    836 => 30,
    837 => 30,
    838 => 30,
    839 => 30,
    840 => 30,
    841 => 30,
    842 => 30,
    843 => 30,
    844 => 30,
    845 => 30,
    846 => 30,
    847 => 30,
    848 => 30,
    849 => 30,
    850 => 30,
    851 => 30,
    852 => 30,
    853 => 30,
    854 => 30,
    855 => 30,
    856 => 30,
    857 => 30,
    858 => 30,
    859 => 30,
    860 => 30,
    861 => 30,
    862 => 30,
    863 => 30,
    864 => 30,
    865 => 30,
    866 => 30,
    867 => 30,
    868 => 30,
    869 => 30,
    870 => 30,
    871 => 30,
    872 => 30,
    873 => 30,
    874 => 30,
    875 => 30,
    876 => 30,
    877 => 30,
    878 => 30,
    879 => 30,
    880 => 30,
    881 => 30,
    882 => 30,
    883 => 30,
    884 => 30,
    885 => 30,
    886 => 30,
    887 => 30,
    888 => 30,
    889 => 30,
    890 => 30,
    891 => 30,
    892 => 30,
    893 => 30,
    894 => 30,
    895 => 30,
    896 => 30,
    897 => 30,
    898 => 30,
    899 => 30,
    900 => 30,
    901 => 30,
    902 => 30,
    903 => 30,
    904 => 30,
    905 => 30,
    906 => 30,
    907 => 31,
    908 => 31,
    909 => 31,
    910 => 31,
    911 => 31,
    912 => 31,
    913 => 31,
    914 => 31,
    915 => 31,
    916 => 31,
    917 => 31,
    918 => 31,
    919 => 31,
    920 => 31,
    921 => 31,
    922 => 31,
    923 => 31,
    924 => 31,
    925 => 31,
    926 => 31,
    927 => 31,
    928 => 31,
    929 => 31,
    930 => 31,
    931 => 31,
    932 => 31,
    933 => 31,
    934 => 31,
    935 => 31,
    936 => 31,
    937 => 31,
    938 => 31,
    939 => 31,
    940 => 31,
    941 => 31,
    942 => 31,
    943 => 31,
    944 => 31,
    945 => 31,
    946 => 31,
    947 => 31,
    948 => 31,
    949 => 31,
    950 => 31,
    951 => 31,
    952 => 31,
    953 => 31,
    954 => 31,
    955 => 31,
    956 => 31,
    957 => 31,
    958 => 31,
    959 => 31,
    960 => 31,
    961 => 31,
    962 => 31,
    963 => 31,
    964 => 31,
    965 => 31,
    966 => 31,
    967 => 31,
    968 => 31,
    969 => 31,
    970 => 31,
    971 => 31,
    972 => 31,
    973 => 31,
    974 => 31,
    975 => 31,
    976 => 31,
    977 => 31,
    978 => 31,
    979 => 31,
    980 => 31,
    981 => 31,
    982 => 31,
    983 => 31,
    984 => 31,
    985 => 31,
    986 => 31,
    987 => 31,
    988 => 31,
    989 => 31,
    990 => 31,
    991 => 31,
    992 => 31,
    993 => 31,
    994 => 31,
    995 => 31,
    996 => 31,
    997 => 31,
    998 => 31,
    999 => 31,
    1000 => 31,
    1001 => 31,
    1002 => 31,
    1003 => 31,
    1004 => 31,
    1005 => 31,
    1006 => 31,
    1007 => 31,
    1008 => 31,
    1009 => 31,
    1010 => 31,
    1011 => 31,
    1012 => 31,
    1013 => 31,
    1014 => 31,
    1015 => 31,
    1016 => 31,
    1017 => 31,
    1018 => 31,
    1019 => 31,
    1020 => 31,
    1021 => 31,
    1022 => 31,
    1023 => 31
  );

begin
  ddfs_out <= std_logic_vector(to_signed(LUT(to_integer(unsigned(address))),6));
end architecture;
